-- NIOSIImicro.vhd

-- Generated using ACDS version 13.0sp1 232 at 2014.10.21.11:37:22

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity NIOSIImicro is
	port (
		clk_50_clk               : in    std_logic                     := '0';             --            clk_50.clk
		sdram_controller_addr    : out   std_logic_vector(11 downto 0);                    --  sdram_controller.addr
		sdram_controller_ba      : out   std_logic_vector(1 downto 0);                     --                  .ba
		sdram_controller_cas_n   : out   std_logic;                                        --                  .cas_n
		sdram_controller_cke     : out   std_logic;                                        --                  .cke
		sdram_controller_cs_n    : out   std_logic;                                        --                  .cs_n
		sdram_controller_dq      : inout std_logic_vector(15 downto 0) := (others => '0'); --                  .dq
		sdram_controller_dqm     : out   std_logic_vector(1 downto 0);                     --                  .dqm
		sdram_controller_ras_n   : out   std_logic;                                        --                  .ras_n
		sdram_controller_we_n    : out   std_logic;                                        --                  .we_n
		pio_in_sw_export         : in    std_logic_vector(17 downto 0) := (others => '0'); --         pio_in_sw.export
		pio_in_key_edge_export   : in    std_logic_vector(2 downto 0)  := (others => '0'); --   pio_in_key_edge.export
		pio_in_ext_export        : in    std_logic_vector(7 downto 0)  := (others => '0'); --        pio_in_ext.export
		pio_out_red_export       : out   std_logic_vector(17 downto 0);                    --       pio_out_red.export
		pio_out_green_export     : out   std_logic_vector(8 downto 0);                     --     pio_out_green.export
		pio_out_ext_export       : out   std_logic_vector(7 downto 0);                     --       pio_out_ext.export
		pio_en_mux_export        : out   std_logic;                                        --        pio_en_mux.export
		pio_direc_export         : out   std_logic_vector(3 downto 0);                     --         pio_direc.export
		pio_direc_ram_export     : out   std_logic_vector(5 downto 0);                     --     pio_direc_ram.export
		pio_wr_export            : out   std_logic;                                        --            pio_wr.export
		pio_sel_salida_export    : out   std_logic_vector(3 downto 0);                     --    pio_sel_salida.export
		pio_datos_export         : out   std_logic_vector(31 downto 0);                    --         pio_datos.export
		pio_compara_int_0_export : in    std_logic                     := '0';             -- pio_compara_int_0.export
		pio_compara_int_1_export : in    std_logic                     := '0';             -- pio_compara_int_1.export
		pio_compara_int_2_export : in    std_logic                     := '0';             -- pio_compara_int_2.export
		pio_compara_int_3_export : in    std_logic                     := '0';             -- pio_compara_int_3.export
		pio_compara_int_4_export : in    std_logic                     := '0';             -- pio_compara_int_4.export
		pio_captura_0_export     : in    std_logic                     := '0';             --     pio_captura_0.export
		pio_captura_1_export     : in    std_logic                     := '0';             --     pio_captura_1.export
		pio_captura_2_export     : in    std_logic                     := '0';             --     pio_captura_2.export
		pio_captura_3_export     : in    std_logic                     := '0';             --     pio_captura_3.export
		pio_captura_4_export     : in    std_logic                     := '0';             --     pio_captura_4.export
		pio_in_32_export         : in    std_logic_vector(31 downto 0) := (others => '0'); --         pio_in_32.export
		lcd_RS                   : out   std_logic;                                        --               lcd.RS
		lcd_RW                   : out   std_logic;                                        --                  .RW
		lcd_data                 : inout std_logic_vector(7 downto 0)  := (others => '0'); --                  .data
		lcd_E                    : out   std_logic;                                        --                  .E
		dm9000a_iOSC_50          : in    std_logic                     := '0';             --           dm9000a.iOSC_50
		dm9000a_ENET_DATA        : inout std_logic_vector(15 downto 0) := (others => '0'); --                  .ENET_DATA
		dm9000a_ENET_CMD         : out   std_logic;                                        --                  .ENET_CMD
		dm9000a_ENET_RD_N        : out   std_logic;                                        --                  .ENET_RD_N
		dm9000a_ENET_WR_N        : out   std_logic;                                        --                  .ENET_WR_N
		dm9000a_ENET_CS_N        : out   std_logic;                                        --                  .ENET_CS_N
		dm9000a_ENET_RST_N       : out   std_logic;                                        --                  .ENET_RST_N
		dm9000a_ENET_CLK         : out   std_logic;                                        --                  .ENET_CLK
		dm9000a_ENET_INT         : in    std_logic                     := '0';             --                  .ENET_INT
		pio_async_reset_export   : out   std_logic;                                        --   pio_async_reset.export
		reset_reset_n            : in    std_logic                     := '0';             --             reset.reset_n
		clock_100_clk            : out   std_logic;                                        --         clock_100.clk
		sdram_clock_clk          : out   std_logic                                         --       sdram_clock.clk
	);
end entity NIOSIImicro;

architecture rtl of NIOSIImicro is
	component NIOSIImicro_cpu is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(24 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(24 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component NIOSIImicro_cpu;

	component NIOSIImicro_pll is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X';             -- write
			address   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0        : out std_logic;                                        -- clk
			c1        : out std_logic;                                        -- clk
			c2        : out std_logic;                                        -- clk
			areset    : in  std_logic                     := 'X';             -- export
			locked    : out std_logic;                                        -- export
			phasedone : out std_logic                                         -- export
		);
	end component NIOSIImicro_pll;

	component NIOSIImicro_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component NIOSIImicro_sdram;

	component NIOSIImicro_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component NIOSIImicro_uart;

	component NIOSIImicro_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component NIOSIImicro_timer_0;

	component NIOSIImicro_timer_1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component NIOSIImicro_timer_1;

	component NIOSIImicro_pio_in_sw is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(17 downto 0) := (others => 'X')  -- export
		);
	end component NIOSIImicro_pio_in_sw;

	component NIOSIImicro_pio_in_key_edge is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component NIOSIImicro_pio_in_key_edge;

	component NIOSIImicro_pio_in_ext is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component NIOSIImicro_pio_in_ext;

	component NIOSIImicro_pio_out_red is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(17 downto 0)                     -- export
		);
	end component NIOSIImicro_pio_out_red;

	component NIOSIImicro_pio_out_green is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(8 downto 0)                      -- export
		);
	end component NIOSIImicro_pio_out_green;

	component NIOSIImicro_pio_out_ext is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component NIOSIImicro_pio_out_ext;

	component NIOSIImicro_pio_en_mux is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component NIOSIImicro_pio_en_mux;

	component NIOSIImicro_pio_direc is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component NIOSIImicro_pio_direc;

	component NIOSIImicro_pio_direc_ram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(5 downto 0)                      -- export
		);
	end component NIOSIImicro_pio_direc_ram;

	component NIOSIImicro_pio_datos is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component NIOSIImicro_pio_datos;

	component NIOSIImicro_pio_compara_int_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component NIOSIImicro_pio_compara_int_0;

	component NIOSIImicro_pio_in_32 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component NIOSIImicro_pio_in_32;

	component NIOSIImicro_lcd is
		port (
			reset_n       : in    std_logic                    := 'X';             -- reset_n
			clk           : in    std_logic                    := 'X';             -- clk
			begintransfer : in    std_logic                    := 'X';             -- begintransfer
			read          : in    std_logic                    := 'X';             -- read
			write         : in    std_logic                    := 'X';             -- write
			readdata      : out   std_logic_vector(7 downto 0);                    -- readdata
			writedata     : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			address       : in    std_logic_vector(1 downto 0) := (others => 'X'); -- address
			LCD_RS        : out   std_logic;                                       -- export
			LCD_RW        : out   std_logic;                                       -- export
			LCD_data      : inout std_logic_vector(7 downto 0) := (others => 'X'); -- export
			LCD_E         : out   std_logic                                        -- export
		);
	end component NIOSIImicro_lcd;

	component NIOSIImicro_system_id is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component NIOSIImicro_system_id;

	component DM9000A_IF is
		port (
			iCLK       : in    std_logic                     := 'X';             -- clk
			iRST_N     : in    std_logic                     := 'X';             -- reset_n
			iOSC_50    : in    std_logic                     := 'X';             -- export
			ENET_DATA  : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			ENET_CMD   : out   std_logic;                                        -- export
			ENET_RD_N  : out   std_logic;                                        -- export
			ENET_WR_N  : out   std_logic;                                        -- export
			ENET_CS_N  : out   std_logic;                                        -- export
			ENET_RST_N : out   std_logic;                                        -- export
			ENET_CLK   : out   std_logic;                                        -- export
			ENET_INT   : in    std_logic                     := 'X';             -- export
			iDATA      : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			iCMD       : in    std_logic                     := 'X';             -- address
			iRD_N      : in    std_logic                     := 'X';             -- read_n
			iWR_N      : in    std_logic                     := 'X';             -- write_n
			iCS_N      : in    std_logic                     := 'X';             -- chipselect_n
			oDATA      : out   std_logic_vector(15 downto 0);                    -- readdata
			oINT       : out   std_logic                                         -- irq
		);
	end component DM9000A_IF;

	component altera_merlin_master_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			av_address              : in  std_logic_vector(24 downto 0)  := (others => 'X'); -- address
			av_write                : in  std_logic                      := 'X';             -- write
			av_read                 : in  std_logic                      := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                     -- readdata
			av_waitrequest          : out std_logic;                                         -- waitrequest
			av_readdatavalid        : out std_logic;                                         -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                      := 'X';             -- debugaccess
			av_lock                 : in  std_logic                      := 'X';             -- lock
			cp_valid                : out std_logic;                                         -- valid
			cp_data                 : out std_logic_vector(103 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_endofpacket          : out std_logic;                                         -- endofpacket
			cp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : in  std_logic                      := 'X';             -- valid
			rp_data                 : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                         -- ready
			av_response             : out std_logic_vector(1 downto 0);                      -- response
			av_writeresponserequest : in  std_logic                      := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                          -- writeresponsevalid
		);
	end component altera_merlin_master_agent;

	component NIOSIImicro_addr_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(103 downto 0);                    -- data
			src_channel        : out std_logic_vector(32 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component NIOSIImicro_addr_router;

	component NIOSIImicro_addr_router_001 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(103 downto 0);                    -- data
			src_channel        : out std_logic_vector(32 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component NIOSIImicro_addr_router_001;

	component NIOSIImicro_id_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(103 downto 0);                    -- data
			src_channel        : out std_logic_vector(32 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component NIOSIImicro_id_router;

	component NIOSIImicro_id_router_001 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(85 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(85 downto 0);                    -- data
			src_channel        : out std_logic_vector(32 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component NIOSIImicro_id_router_001;

	component NIOSIImicro_id_router_003 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(103 downto 0);                    -- data
			src_channel        : out std_logic_vector(32 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component NIOSIImicro_id_router_003;

	component altera_merlin_traffic_limiter is
		generic (
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_TRANS_POSTED          : integer := 0;
			PKT_TRANS_WRITE           : integer := 0;
			MAX_OUTSTANDING_RESPONSES : integer := 0;
			PIPELINED                 : integer := 0;
			ST_DATA_W                 : integer := 72;
			ST_CHANNEL_W              : integer := 1;
			VALID_WIDTH               : integer := 1;
			ENFORCE_ORDER             : integer := 1;
			PREVENT_HAZARDS           : integer := 0;
			PKT_BYTE_CNT_H            : integer := 0;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 0;
			PKT_BYTEEN_L              : integer := 0
		);
		port (
			clk                    : in  std_logic                      := 'X';             -- clk
			reset                  : in  std_logic                      := 'X';             -- reset
			cmd_sink_ready         : out std_logic;                                         -- ready
			cmd_sink_valid         : in  std_logic                      := 'X';             -- valid
			cmd_sink_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			cmd_sink_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			cmd_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			cmd_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			cmd_src_ready          : in  std_logic                      := 'X';             -- ready
			cmd_src_data           : out std_logic_vector(103 downto 0);                    -- data
			cmd_src_channel        : out std_logic_vector(32 downto 0);                     -- channel
			cmd_src_startofpacket  : out std_logic;                                         -- startofpacket
			cmd_src_endofpacket    : out std_logic;                                         -- endofpacket
			rsp_sink_ready         : out std_logic;                                         -- ready
			rsp_sink_valid         : in  std_logic                      := 'X';             -- valid
			rsp_sink_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			rsp_sink_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			rsp_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			rsp_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			rsp_src_ready          : in  std_logic                      := 'X';             -- ready
			rsp_src_valid          : out std_logic;                                         -- valid
			rsp_src_data           : out std_logic_vector(103 downto 0);                    -- data
			rsp_src_channel        : out std_logic_vector(32 downto 0);                     -- channel
			rsp_src_startofpacket  : out std_logic;                                         -- startofpacket
			rsp_src_endofpacket    : out std_logic;                                         -- endofpacket
			cmd_src_valid          : out std_logic_vector(32 downto 0)                      -- data
		);
	end component altera_merlin_traffic_limiter;

	component altera_merlin_burst_adapter is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			sink0_valid           : in  std_logic                     := 'X';             -- valid
			sink0_data            : in  std_logic_vector(85 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(32 downto 0) := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                        -- ready
			source0_valid         : out std_logic;                                        -- valid
			source0_data          : out std_logic_vector(85 downto 0);                    -- data
			source0_channel       : out std_logic_vector(32 downto 0);                    -- channel
			source0_startofpacket : out std_logic;                                        -- startofpacket
			source0_endofpacket   : out std_logic;                                        -- endofpacket
			source0_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component altera_merlin_burst_adapter;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component altera_reset_controller;

	component NIOSIImicro_cmd_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- data
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(103 downto 0);                    -- data
			src0_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(103 downto 0);                    -- data
			src1_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic;                                         -- endofpacket
			src2_ready         : in  std_logic                      := 'X';             -- ready
			src2_valid         : out std_logic;                                         -- valid
			src2_data          : out std_logic_vector(103 downto 0);                    -- data
			src2_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src2_startofpacket : out std_logic;                                         -- startofpacket
			src2_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component NIOSIImicro_cmd_xbar_demux;

	component NIOSIImicro_cmd_xbar_demux_001 is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			sink_ready          : out std_logic;                                         -- ready
			sink_channel        : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink_data           : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink_valid          : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready          : in  std_logic                      := 'X';             -- ready
			src0_valid          : out std_logic;                                         -- valid
			src0_data           : out std_logic_vector(103 downto 0);                    -- data
			src0_channel        : out std_logic_vector(32 downto 0);                     -- channel
			src0_startofpacket  : out std_logic;                                         -- startofpacket
			src0_endofpacket    : out std_logic;                                         -- endofpacket
			src1_ready          : in  std_logic                      := 'X';             -- ready
			src1_valid          : out std_logic;                                         -- valid
			src1_data           : out std_logic_vector(103 downto 0);                    -- data
			src1_channel        : out std_logic_vector(32 downto 0);                     -- channel
			src1_startofpacket  : out std_logic;                                         -- startofpacket
			src1_endofpacket    : out std_logic;                                         -- endofpacket
			src2_ready          : in  std_logic                      := 'X';             -- ready
			src2_valid          : out std_logic;                                         -- valid
			src2_data           : out std_logic_vector(103 downto 0);                    -- data
			src2_channel        : out std_logic_vector(32 downto 0);                     -- channel
			src2_startofpacket  : out std_logic;                                         -- startofpacket
			src2_endofpacket    : out std_logic;                                         -- endofpacket
			src3_ready          : in  std_logic                      := 'X';             -- ready
			src3_valid          : out std_logic;                                         -- valid
			src3_data           : out std_logic_vector(103 downto 0);                    -- data
			src3_channel        : out std_logic_vector(32 downto 0);                     -- channel
			src3_startofpacket  : out std_logic;                                         -- startofpacket
			src3_endofpacket    : out std_logic;                                         -- endofpacket
			src4_ready          : in  std_logic                      := 'X';             -- ready
			src4_valid          : out std_logic;                                         -- valid
			src4_data           : out std_logic_vector(103 downto 0);                    -- data
			src4_channel        : out std_logic_vector(32 downto 0);                     -- channel
			src4_startofpacket  : out std_logic;                                         -- startofpacket
			src4_endofpacket    : out std_logic;                                         -- endofpacket
			src5_ready          : in  std_logic                      := 'X';             -- ready
			src5_valid          : out std_logic;                                         -- valid
			src5_data           : out std_logic_vector(103 downto 0);                    -- data
			src5_channel        : out std_logic_vector(32 downto 0);                     -- channel
			src5_startofpacket  : out std_logic;                                         -- startofpacket
			src5_endofpacket    : out std_logic;                                         -- endofpacket
			src6_ready          : in  std_logic                      := 'X';             -- ready
			src6_valid          : out std_logic;                                         -- valid
			src6_data           : out std_logic_vector(103 downto 0);                    -- data
			src6_channel        : out std_logic_vector(32 downto 0);                     -- channel
			src6_startofpacket  : out std_logic;                                         -- startofpacket
			src6_endofpacket    : out std_logic;                                         -- endofpacket
			src7_ready          : in  std_logic                      := 'X';             -- ready
			src7_valid          : out std_logic;                                         -- valid
			src7_data           : out std_logic_vector(103 downto 0);                    -- data
			src7_channel        : out std_logic_vector(32 downto 0);                     -- channel
			src7_startofpacket  : out std_logic;                                         -- startofpacket
			src7_endofpacket    : out std_logic;                                         -- endofpacket
			src8_ready          : in  std_logic                      := 'X';             -- ready
			src8_valid          : out std_logic;                                         -- valid
			src8_data           : out std_logic_vector(103 downto 0);                    -- data
			src8_channel        : out std_logic_vector(32 downto 0);                     -- channel
			src8_startofpacket  : out std_logic;                                         -- startofpacket
			src8_endofpacket    : out std_logic;                                         -- endofpacket
			src9_ready          : in  std_logic                      := 'X';             -- ready
			src9_valid          : out std_logic;                                         -- valid
			src9_data           : out std_logic_vector(103 downto 0);                    -- data
			src9_channel        : out std_logic_vector(32 downto 0);                     -- channel
			src9_startofpacket  : out std_logic;                                         -- startofpacket
			src9_endofpacket    : out std_logic;                                         -- endofpacket
			src10_ready         : in  std_logic                      := 'X';             -- ready
			src10_valid         : out std_logic;                                         -- valid
			src10_data          : out std_logic_vector(103 downto 0);                    -- data
			src10_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src10_startofpacket : out std_logic;                                         -- startofpacket
			src10_endofpacket   : out std_logic;                                         -- endofpacket
			src11_ready         : in  std_logic                      := 'X';             -- ready
			src11_valid         : out std_logic;                                         -- valid
			src11_data          : out std_logic_vector(103 downto 0);                    -- data
			src11_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src11_startofpacket : out std_logic;                                         -- startofpacket
			src11_endofpacket   : out std_logic;                                         -- endofpacket
			src12_ready         : in  std_logic                      := 'X';             -- ready
			src12_valid         : out std_logic;                                         -- valid
			src12_data          : out std_logic_vector(103 downto 0);                    -- data
			src12_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src12_startofpacket : out std_logic;                                         -- startofpacket
			src12_endofpacket   : out std_logic;                                         -- endofpacket
			src13_ready         : in  std_logic                      := 'X';             -- ready
			src13_valid         : out std_logic;                                         -- valid
			src13_data          : out std_logic_vector(103 downto 0);                    -- data
			src13_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src13_startofpacket : out std_logic;                                         -- startofpacket
			src13_endofpacket   : out std_logic;                                         -- endofpacket
			src14_ready         : in  std_logic                      := 'X';             -- ready
			src14_valid         : out std_logic;                                         -- valid
			src14_data          : out std_logic_vector(103 downto 0);                    -- data
			src14_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src14_startofpacket : out std_logic;                                         -- startofpacket
			src14_endofpacket   : out std_logic;                                         -- endofpacket
			src15_ready         : in  std_logic                      := 'X';             -- ready
			src15_valid         : out std_logic;                                         -- valid
			src15_data          : out std_logic_vector(103 downto 0);                    -- data
			src15_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src15_startofpacket : out std_logic;                                         -- startofpacket
			src15_endofpacket   : out std_logic;                                         -- endofpacket
			src16_ready         : in  std_logic                      := 'X';             -- ready
			src16_valid         : out std_logic;                                         -- valid
			src16_data          : out std_logic_vector(103 downto 0);                    -- data
			src16_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src16_startofpacket : out std_logic;                                         -- startofpacket
			src16_endofpacket   : out std_logic;                                         -- endofpacket
			src17_ready         : in  std_logic                      := 'X';             -- ready
			src17_valid         : out std_logic;                                         -- valid
			src17_data          : out std_logic_vector(103 downto 0);                    -- data
			src17_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src17_startofpacket : out std_logic;                                         -- startofpacket
			src17_endofpacket   : out std_logic;                                         -- endofpacket
			src18_ready         : in  std_logic                      := 'X';             -- ready
			src18_valid         : out std_logic;                                         -- valid
			src18_data          : out std_logic_vector(103 downto 0);                    -- data
			src18_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src18_startofpacket : out std_logic;                                         -- startofpacket
			src18_endofpacket   : out std_logic;                                         -- endofpacket
			src19_ready         : in  std_logic                      := 'X';             -- ready
			src19_valid         : out std_logic;                                         -- valid
			src19_data          : out std_logic_vector(103 downto 0);                    -- data
			src19_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src19_startofpacket : out std_logic;                                         -- startofpacket
			src19_endofpacket   : out std_logic;                                         -- endofpacket
			src20_ready         : in  std_logic                      := 'X';             -- ready
			src20_valid         : out std_logic;                                         -- valid
			src20_data          : out std_logic_vector(103 downto 0);                    -- data
			src20_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src20_startofpacket : out std_logic;                                         -- startofpacket
			src20_endofpacket   : out std_logic;                                         -- endofpacket
			src21_ready         : in  std_logic                      := 'X';             -- ready
			src21_valid         : out std_logic;                                         -- valid
			src21_data          : out std_logic_vector(103 downto 0);                    -- data
			src21_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src21_startofpacket : out std_logic;                                         -- startofpacket
			src21_endofpacket   : out std_logic;                                         -- endofpacket
			src22_ready         : in  std_logic                      := 'X';             -- ready
			src22_valid         : out std_logic;                                         -- valid
			src22_data          : out std_logic_vector(103 downto 0);                    -- data
			src22_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src22_startofpacket : out std_logic;                                         -- startofpacket
			src22_endofpacket   : out std_logic;                                         -- endofpacket
			src23_ready         : in  std_logic                      := 'X';             -- ready
			src23_valid         : out std_logic;                                         -- valid
			src23_data          : out std_logic_vector(103 downto 0);                    -- data
			src23_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src23_startofpacket : out std_logic;                                         -- startofpacket
			src23_endofpacket   : out std_logic;                                         -- endofpacket
			src24_ready         : in  std_logic                      := 'X';             -- ready
			src24_valid         : out std_logic;                                         -- valid
			src24_data          : out std_logic_vector(103 downto 0);                    -- data
			src24_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src24_startofpacket : out std_logic;                                         -- startofpacket
			src24_endofpacket   : out std_logic;                                         -- endofpacket
			src25_ready         : in  std_logic                      := 'X';             -- ready
			src25_valid         : out std_logic;                                         -- valid
			src25_data          : out std_logic_vector(103 downto 0);                    -- data
			src25_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src25_startofpacket : out std_logic;                                         -- startofpacket
			src25_endofpacket   : out std_logic;                                         -- endofpacket
			src26_ready         : in  std_logic                      := 'X';             -- ready
			src26_valid         : out std_logic;                                         -- valid
			src26_data          : out std_logic_vector(103 downto 0);                    -- data
			src26_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src26_startofpacket : out std_logic;                                         -- startofpacket
			src26_endofpacket   : out std_logic;                                         -- endofpacket
			src27_ready         : in  std_logic                      := 'X';             -- ready
			src27_valid         : out std_logic;                                         -- valid
			src27_data          : out std_logic_vector(103 downto 0);                    -- data
			src27_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src27_startofpacket : out std_logic;                                         -- startofpacket
			src27_endofpacket   : out std_logic;                                         -- endofpacket
			src28_ready         : in  std_logic                      := 'X';             -- ready
			src28_valid         : out std_logic;                                         -- valid
			src28_data          : out std_logic_vector(103 downto 0);                    -- data
			src28_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src28_startofpacket : out std_logic;                                         -- startofpacket
			src28_endofpacket   : out std_logic;                                         -- endofpacket
			src29_ready         : in  std_logic                      := 'X';             -- ready
			src29_valid         : out std_logic;                                         -- valid
			src29_data          : out std_logic_vector(103 downto 0);                    -- data
			src29_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src29_startofpacket : out std_logic;                                         -- startofpacket
			src29_endofpacket   : out std_logic;                                         -- endofpacket
			src30_ready         : in  std_logic                      := 'X';             -- ready
			src30_valid         : out std_logic;                                         -- valid
			src30_data          : out std_logic_vector(103 downto 0);                    -- data
			src30_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src30_startofpacket : out std_logic;                                         -- startofpacket
			src30_endofpacket   : out std_logic;                                         -- endofpacket
			src31_ready         : in  std_logic                      := 'X';             -- ready
			src31_valid         : out std_logic;                                         -- valid
			src31_data          : out std_logic_vector(103 downto 0);                    -- data
			src31_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src31_startofpacket : out std_logic;                                         -- startofpacket
			src31_endofpacket   : out std_logic;                                         -- endofpacket
			src32_ready         : in  std_logic                      := 'X';             -- ready
			src32_valid         : out std_logic;                                         -- valid
			src32_data          : out std_logic_vector(103 downto 0);                    -- data
			src32_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src32_startofpacket : out std_logic;                                         -- startofpacket
			src32_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component NIOSIImicro_cmd_xbar_demux_001;

	component NIOSIImicro_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(103 downto 0);                    -- data
			src_channel         : out std_logic_vector(32 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component NIOSIImicro_cmd_xbar_mux;

	component NIOSIImicro_rsp_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(103 downto 0);                    -- data
			src0_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(103 downto 0);                    -- data
			src1_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component NIOSIImicro_rsp_xbar_demux;

	component NIOSIImicro_rsp_xbar_demux_003 is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(103 downto 0);                    -- data
			src0_channel       : out std_logic_vector(32 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component NIOSIImicro_rsp_xbar_demux_003;

	component NIOSIImicro_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(103 downto 0);                    -- data
			src_channel         : out std_logic_vector(32 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                         -- ready
			sink2_valid         : in  std_logic                      := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component NIOSIImicro_rsp_xbar_mux;

	component NIOSIImicro_rsp_xbar_mux_001 is
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			src_ready            : in  std_logic                      := 'X';             -- ready
			src_valid            : out std_logic;                                         -- valid
			src_data             : out std_logic_vector(103 downto 0);                    -- data
			src_channel          : out std_logic_vector(32 downto 0);                     -- channel
			src_startofpacket    : out std_logic;                                         -- startofpacket
			src_endofpacket      : out std_logic;                                         -- endofpacket
			sink0_ready          : out std_logic;                                         -- ready
			sink0_valid          : in  std_logic                      := 'X';             -- valid
			sink0_channel        : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink0_data           : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink0_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready          : out std_logic;                                         -- ready
			sink1_valid          : in  std_logic                      := 'X';             -- valid
			sink1_channel        : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink1_data           : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink1_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink2_ready          : out std_logic;                                         -- ready
			sink2_valid          : in  std_logic                      := 'X';             -- valid
			sink2_channel        : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink2_data           : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink2_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink2_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink3_ready          : out std_logic;                                         -- ready
			sink3_valid          : in  std_logic                      := 'X';             -- valid
			sink3_channel        : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink3_data           : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink3_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink3_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink4_ready          : out std_logic;                                         -- ready
			sink4_valid          : in  std_logic                      := 'X';             -- valid
			sink4_channel        : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink4_data           : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink4_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink4_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink5_ready          : out std_logic;                                         -- ready
			sink5_valid          : in  std_logic                      := 'X';             -- valid
			sink5_channel        : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink5_data           : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink5_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink5_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink6_ready          : out std_logic;                                         -- ready
			sink6_valid          : in  std_logic                      := 'X';             -- valid
			sink6_channel        : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink6_data           : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink6_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink6_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink7_ready          : out std_logic;                                         -- ready
			sink7_valid          : in  std_logic                      := 'X';             -- valid
			sink7_channel        : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink7_data           : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink7_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink7_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink8_ready          : out std_logic;                                         -- ready
			sink8_valid          : in  std_logic                      := 'X';             -- valid
			sink8_channel        : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink8_data           : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink8_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink8_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink9_ready          : out std_logic;                                         -- ready
			sink9_valid          : in  std_logic                      := 'X';             -- valid
			sink9_channel        : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink9_data           : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink9_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink9_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink10_ready         : out std_logic;                                         -- ready
			sink10_valid         : in  std_logic                      := 'X';             -- valid
			sink10_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink10_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink10_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink10_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink11_ready         : out std_logic;                                         -- ready
			sink11_valid         : in  std_logic                      := 'X';             -- valid
			sink11_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink11_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink11_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink11_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink12_ready         : out std_logic;                                         -- ready
			sink12_valid         : in  std_logic                      := 'X';             -- valid
			sink12_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink12_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink12_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink12_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink13_ready         : out std_logic;                                         -- ready
			sink13_valid         : in  std_logic                      := 'X';             -- valid
			sink13_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink13_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink13_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink13_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink14_ready         : out std_logic;                                         -- ready
			sink14_valid         : in  std_logic                      := 'X';             -- valid
			sink14_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink14_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink14_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink14_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink15_ready         : out std_logic;                                         -- ready
			sink15_valid         : in  std_logic                      := 'X';             -- valid
			sink15_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink15_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink15_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink15_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink16_ready         : out std_logic;                                         -- ready
			sink16_valid         : in  std_logic                      := 'X';             -- valid
			sink16_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink16_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink16_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink16_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink17_ready         : out std_logic;                                         -- ready
			sink17_valid         : in  std_logic                      := 'X';             -- valid
			sink17_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink17_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink17_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink17_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink18_ready         : out std_logic;                                         -- ready
			sink18_valid         : in  std_logic                      := 'X';             -- valid
			sink18_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink18_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink18_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink18_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink19_ready         : out std_logic;                                         -- ready
			sink19_valid         : in  std_logic                      := 'X';             -- valid
			sink19_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink19_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink19_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink19_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink20_ready         : out std_logic;                                         -- ready
			sink20_valid         : in  std_logic                      := 'X';             -- valid
			sink20_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink20_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink20_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink20_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink21_ready         : out std_logic;                                         -- ready
			sink21_valid         : in  std_logic                      := 'X';             -- valid
			sink21_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink21_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink21_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink21_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink22_ready         : out std_logic;                                         -- ready
			sink22_valid         : in  std_logic                      := 'X';             -- valid
			sink22_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink22_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink22_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink22_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink23_ready         : out std_logic;                                         -- ready
			sink23_valid         : in  std_logic                      := 'X';             -- valid
			sink23_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink23_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink23_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink23_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink24_ready         : out std_logic;                                         -- ready
			sink24_valid         : in  std_logic                      := 'X';             -- valid
			sink24_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink24_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink24_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink24_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink25_ready         : out std_logic;                                         -- ready
			sink25_valid         : in  std_logic                      := 'X';             -- valid
			sink25_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink25_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink25_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink25_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink26_ready         : out std_logic;                                         -- ready
			sink26_valid         : in  std_logic                      := 'X';             -- valid
			sink26_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink26_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink26_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink26_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink27_ready         : out std_logic;                                         -- ready
			sink27_valid         : in  std_logic                      := 'X';             -- valid
			sink27_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink27_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink27_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink27_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink28_ready         : out std_logic;                                         -- ready
			sink28_valid         : in  std_logic                      := 'X';             -- valid
			sink28_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink28_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink28_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink28_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink29_ready         : out std_logic;                                         -- ready
			sink29_valid         : in  std_logic                      := 'X';             -- valid
			sink29_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink29_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink29_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink29_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink30_ready         : out std_logic;                                         -- ready
			sink30_valid         : in  std_logic                      := 'X';             -- valid
			sink30_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink30_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink30_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink30_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink31_ready         : out std_logic;                                         -- ready
			sink31_valid         : in  std_logic                      := 'X';             -- valid
			sink31_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink31_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink31_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink31_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink32_ready         : out std_logic;                                         -- ready
			sink32_valid         : in  std_logic                      := 'X';             -- valid
			sink32_channel       : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			sink32_data          : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			sink32_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink32_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component NIOSIImicro_rsp_xbar_mux_001;

	component altera_avalon_st_handshake_clock_crosser is
		generic (
			DATA_WIDTH          : integer := 8;
			BITS_PER_SYMBOL     : integer := 8;
			USE_PACKETS         : integer := 0;
			USE_CHANNEL         : integer := 0;
			CHANNEL_WIDTH       : integer := 1;
			USE_ERROR           : integer := 0;
			ERROR_WIDTH         : integer := 1;
			VALID_SYNC_DEPTH    : integer := 2;
			READY_SYNC_DEPTH    : integer := 2;
			USE_OUTPUT_PIPELINE : integer := 1
		);
		port (
			in_clk            : in  std_logic                      := 'X';             -- clk
			in_reset          : in  std_logic                      := 'X';             -- reset
			out_clk           : in  std_logic                      := 'X';             -- clk
			out_reset         : in  std_logic                      := 'X';             -- reset
			in_ready          : out std_logic;                                         -- ready
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			in_channel        : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			in_data           : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_valid         : out std_logic;                                         -- valid
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			out_channel       : out std_logic_vector(32 downto 0);                     -- channel
			out_data          : out std_logic_vector(103 downto 0);                    -- data
			in_empty          : in  std_logic                      := 'X';             -- empty
			in_error          : in  std_logic                      := 'X';             -- error
			out_empty         : out std_logic;                                         -- empty
			out_error         : out std_logic                                          -- error
		);
	end component altera_avalon_st_handshake_clock_crosser;

	component NIOSIImicro_irq_mapper is
		port (
			clk            : in  std_logic                     := 'X'; -- clk
			reset          : in  std_logic                     := 'X'; -- reset
			receiver0_irq  : in  std_logic                     := 'X'; -- irq
			receiver1_irq  : in  std_logic                     := 'X'; -- irq
			receiver2_irq  : in  std_logic                     := 'X'; -- irq
			receiver3_irq  : in  std_logic                     := 'X'; -- irq
			receiver4_irq  : in  std_logic                     := 'X'; -- irq
			receiver5_irq  : in  std_logic                     := 'X'; -- irq
			receiver6_irq  : in  std_logic                     := 'X'; -- irq
			receiver7_irq  : in  std_logic                     := 'X'; -- irq
			receiver8_irq  : in  std_logic                     := 'X'; -- irq
			receiver9_irq  : in  std_logic                     := 'X'; -- irq
			receiver10_irq : in  std_logic                     := 'X'; -- irq
			receiver11_irq : in  std_logic                     := 'X'; -- irq
			receiver12_irq : in  std_logic                     := 'X'; -- irq
			receiver13_irq : in  std_logic                     := 'X'; -- irq
			receiver14_irq : in  std_logic                     := 'X'; -- irq
			receiver15_irq : in  std_logic                     := 'X'; -- irq
			sender_irq     : out std_logic_vector(31 downto 0)         -- irq
		);
	end component NIOSIImicro_irq_mapper;

	component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(104 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(104 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- address
			csr_read          : in  std_logic                      := 'X';             -- read
			csr_write         : in  std_logic                      := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                         -- data
			almost_empty_data : out std_logic;                                         -- data
			in_empty          : in  std_logic                      := 'X';             -- empty
			out_empty         : out std_logic;                                         -- empty
			in_error          : in  std_logic                      := 'X';             -- error
			out_error         : out std_logic;                                         -- error
			in_channel        : in  std_logic                      := 'X';             -- channel
			out_channel       : out std_logic                                          -- channel
		);
	end component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component niosiimicro_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(86 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component niosiimicro_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component niosiimicro_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(17 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component niosiimicro_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component niosiimicro_pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(33 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(33 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component niosiimicro_pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(103 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(104 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(104 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                         -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                      := 'X'              -- writeresponsevalid
		);
	end component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent;

	component niosiimicro_sdram_s1_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(1 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(85 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(85 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(32 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(86 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(86 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(17 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component niosiimicro_sdram_s1_translator_avalon_universal_slave_0_agent;

	component niosiimicro_width_adapter is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(103 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(85 downto 0);                     -- data
			out_channel          : out std_logic_vector(32 downto 0);                     -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component niosiimicro_width_adapter;

	component niosiimicro_width_adapter_001 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(85 downto 0)  := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(103 downto 0);                    -- data
			out_channel          : out std_logic_vector(32 downto 0);                     -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component niosiimicro_width_adapter_001;

	component niosiimicro_cpu_instruction_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(24 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component niosiimicro_cpu_instruction_master_translator;

	component niosiimicro_cpu_data_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(24 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component niosiimicro_cpu_data_master_translator;

	component niosiimicro_cpu_jtag_debug_module_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(8 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component niosiimicro_cpu_jtag_debug_module_translator;

	component niosiimicro_sdram_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(21 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(1 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_writebyteenable       : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component niosiimicro_sdram_s1_translator;

	component niosiimicro_system_id_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component niosiimicro_system_id_control_slave_translator;

	component niosiimicro_pll_pll_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component niosiimicro_pll_pll_slave_translator;

	component niosiimicro_uart_avalon_jtag_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component niosiimicro_uart_avalon_jtag_slave_translator;

	component niosiimicro_timer_0_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component niosiimicro_timer_0_s1_translator;

	component niosiimicro_pio_in_sw_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component niosiimicro_pio_in_sw_s1_translator;

	component niosiimicro_pio_in_key_edge_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component niosiimicro_pio_in_key_edge_s1_translator;

	component niosiimicro_pio_out_red_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component niosiimicro_pio_out_red_s1_translator;

	component niosiimicro_lcd_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(7 downto 0);                     -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component niosiimicro_lcd_control_slave_translator;

	component niosiimicro_dm9000a_avalon_slave_0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component niosiimicro_dm9000a_avalon_slave_0_translator;

	signal pll_c0_clk                                                                                   : std_logic;                      -- pll:c0 -> [DM9000A:iCLK, DM9000A_avalon_slave_0_translator:clk, DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, addr_router_001:clk, burst_adapter:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_002:clk, cpu:clk, cpu_data_master_translator:clk, cpu_data_master_translator_avalon_universal_master_0_agent:clk, cpu_instruction_master_translator:clk, cpu_instruction_master_translator_avalon_universal_master_0_agent:clk, cpu_jtag_debug_module_translator:clk, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, crosser:in_clk, crosser_001:out_clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_015:clk, id_router_016:clk, id_router_017:clk, id_router_018:clk, id_router_019:clk, id_router_020:clk, id_router_021:clk, id_router_022:clk, id_router_023:clk, id_router_024:clk, id_router_025:clk, id_router_026:clk, id_router_027:clk, id_router_028:clk, id_router_029:clk, id_router_030:clk, id_router_031:clk, id_router_032:clk, irq_mapper:clk, lcd:clk, lcd_control_slave_translator:clk, lcd_control_slave_translator_avalon_universal_slave_0_agent:clk, lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter:clk, pio_async_reset:clk, pio_async_reset_s1_translator:clk, pio_async_reset_s1_translator_avalon_universal_slave_0_agent:clk, pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_captura_0:clk, pio_captura_0_s1_translator:clk, pio_captura_0_s1_translator_avalon_universal_slave_0_agent:clk, pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_captura_1:clk, pio_captura_1_s1_translator:clk, pio_captura_1_s1_translator_avalon_universal_slave_0_agent:clk, pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_captura_2:clk, pio_captura_2_s1_translator:clk, pio_captura_2_s1_translator_avalon_universal_slave_0_agent:clk, pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_captura_3:clk, pio_captura_3_s1_translator:clk, pio_captura_3_s1_translator_avalon_universal_slave_0_agent:clk, pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_captura_4:clk, pio_captura_4_s1_translator:clk, pio_captura_4_s1_translator_avalon_universal_slave_0_agent:clk, pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_compara_int_0:clk, pio_compara_int_0_s1_translator:clk, pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:clk, pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_compara_int_1:clk, pio_compara_int_1_s1_translator:clk, pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:clk, pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_compara_int_2:clk, pio_compara_int_2_s1_translator:clk, pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:clk, pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_compara_int_3:clk, pio_compara_int_3_s1_translator:clk, pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:clk, pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_compara_int_4:clk, pio_compara_int_4_s1_translator:clk, pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:clk, pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_datos:clk, pio_datos_s1_translator:clk, pio_datos_s1_translator_avalon_universal_slave_0_agent:clk, pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_direc:clk, pio_direc_ram:clk, pio_direc_ram_s1_translator:clk, pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:clk, pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_direc_s1_translator:clk, pio_direc_s1_translator_avalon_universal_slave_0_agent:clk, pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_en_mux:clk, pio_en_mux_s1_translator:clk, pio_en_mux_s1_translator_avalon_universal_slave_0_agent:clk, pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_in_32:clk, pio_in_32_s1_translator:clk, pio_in_32_s1_translator_avalon_universal_slave_0_agent:clk, pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_in_ext:clk, pio_in_ext_s1_translator:clk, pio_in_ext_s1_translator_avalon_universal_slave_0_agent:clk, pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_in_key_edge:clk, pio_in_key_edge_s1_translator:clk, pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:clk, pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_in_sw:clk, pio_in_sw_s1_translator:clk, pio_in_sw_s1_translator_avalon_universal_slave_0_agent:clk, pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_out_ext:clk, pio_out_ext_s1_translator:clk, pio_out_ext_s1_translator_avalon_universal_slave_0_agent:clk, pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_out_green:clk, pio_out_green_s1_translator:clk, pio_out_green_s1_translator_avalon_universal_slave_0_agent:clk, pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_out_red:clk, pio_out_red_s1_translator:clk, pio_out_red_s1_translator_avalon_universal_slave_0_agent:clk, pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_sel_salida:clk, pio_sel_salida_s1_translator:clk, pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:clk, pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_wr:clk, pio_wr_s1_translator:clk, pio_wr_s1_translator_avalon_universal_slave_0_agent:clk, pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_015:clk, rsp_xbar_demux_016:clk, rsp_xbar_demux_017:clk, rsp_xbar_demux_018:clk, rsp_xbar_demux_019:clk, rsp_xbar_demux_020:clk, rsp_xbar_demux_021:clk, rsp_xbar_demux_022:clk, rsp_xbar_demux_023:clk, rsp_xbar_demux_024:clk, rsp_xbar_demux_025:clk, rsp_xbar_demux_026:clk, rsp_xbar_demux_027:clk, rsp_xbar_demux_028:clk, rsp_xbar_demux_029:clk, rsp_xbar_demux_030:clk, rsp_xbar_demux_031:clk, rsp_xbar_demux_032:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, sdram:clk, sdram_s1_translator:clk, sdram_s1_translator_avalon_universal_slave_0_agent:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, system_id:clock, system_id_control_slave_translator:clk, system_id_control_slave_translator_avalon_universal_slave_0_agent:clk, system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer_0:clk, timer_0_s1_translator:clk, timer_0_s1_translator_avalon_universal_slave_0_agent:clk, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer_1:clk, timer_1_s1_translator:clk, timer_1_s1_translator_avalon_universal_slave_0_agent:clk, timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, uart:clk, uart_avalon_jtag_slave_translator:clk, uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter:clk, width_adapter_001:clk]
	signal cpu_instruction_master_waitrequest                                                           : std_logic;                      -- cpu_instruction_master_translator:av_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                                               : std_logic_vector(24 downto 0);  -- cpu:i_address -> cpu_instruction_master_translator:av_address
	signal cpu_instruction_master_read                                                                  : std_logic;                      -- cpu:i_read -> cpu_instruction_master_translator:av_read
	signal cpu_instruction_master_readdata                                                              : std_logic_vector(31 downto 0);  -- cpu_instruction_master_translator:av_readdata -> cpu:i_readdata
	signal cpu_instruction_master_readdatavalid                                                         : std_logic;                      -- cpu_instruction_master_translator:av_readdatavalid -> cpu:i_readdatavalid
	signal cpu_data_master_waitrequest                                                                  : std_logic;                      -- cpu_data_master_translator:av_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_writedata                                                                    : std_logic_vector(31 downto 0);  -- cpu:d_writedata -> cpu_data_master_translator:av_writedata
	signal cpu_data_master_address                                                                      : std_logic_vector(24 downto 0);  -- cpu:d_address -> cpu_data_master_translator:av_address
	signal cpu_data_master_write                                                                        : std_logic;                      -- cpu:d_write -> cpu_data_master_translator:av_write
	signal cpu_data_master_read                                                                         : std_logic;                      -- cpu:d_read -> cpu_data_master_translator:av_read
	signal cpu_data_master_readdata                                                                     : std_logic_vector(31 downto 0);  -- cpu_data_master_translator:av_readdata -> cpu:d_readdata
	signal cpu_data_master_debugaccess                                                                  : std_logic;                      -- cpu:jtag_debug_module_debugaccess_to_roms -> cpu_data_master_translator:av_debugaccess
	signal cpu_data_master_byteenable                                                                   : std_logic_vector(3 downto 0);   -- cpu:d_byteenable -> cpu_data_master_translator:av_byteenable
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest                             : std_logic;                      -- cpu:jtag_debug_module_waitrequest -> cpu_jtag_debug_module_translator:av_waitrequest
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata                               : std_logic_vector(31 downto 0);  -- cpu_jtag_debug_module_translator:av_writedata -> cpu:jtag_debug_module_writedata
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_address                                 : std_logic_vector(8 downto 0);   -- cpu_jtag_debug_module_translator:av_address -> cpu:jtag_debug_module_address
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_write                                   : std_logic;                      -- cpu_jtag_debug_module_translator:av_write -> cpu:jtag_debug_module_write
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_read                                    : std_logic;                      -- cpu_jtag_debug_module_translator:av_read -> cpu:jtag_debug_module_read
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata                                : std_logic_vector(31 downto 0);  -- cpu:jtag_debug_module_readdata -> cpu_jtag_debug_module_translator:av_readdata
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                             : std_logic;                      -- cpu_jtag_debug_module_translator:av_debugaccess -> cpu:jtag_debug_module_debugaccess
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                              : std_logic_vector(3 downto 0);   -- cpu_jtag_debug_module_translator:av_byteenable -> cpu:jtag_debug_module_byteenable
	signal sdram_s1_translator_avalon_anti_slave_0_waitrequest                                          : std_logic;                      -- sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	signal sdram_s1_translator_avalon_anti_slave_0_writedata                                            : std_logic_vector(15 downto 0);  -- sdram_s1_translator:av_writedata -> sdram:az_data
	signal sdram_s1_translator_avalon_anti_slave_0_address                                              : std_logic_vector(21 downto 0);  -- sdram_s1_translator:av_address -> sdram:az_addr
	signal sdram_s1_translator_avalon_anti_slave_0_chipselect                                           : std_logic;                      -- sdram_s1_translator:av_chipselect -> sdram:az_cs
	signal sdram_s1_translator_avalon_anti_slave_0_write                                                : std_logic;                      -- sdram_s1_translator:av_write -> sdram_s1_translator_avalon_anti_slave_0_write:in
	signal sdram_s1_translator_avalon_anti_slave_0_read                                                 : std_logic;                      -- sdram_s1_translator:av_read -> sdram_s1_translator_avalon_anti_slave_0_read:in
	signal sdram_s1_translator_avalon_anti_slave_0_readdata                                             : std_logic_vector(15 downto 0);  -- sdram:za_data -> sdram_s1_translator:av_readdata
	signal sdram_s1_translator_avalon_anti_slave_0_readdatavalid                                        : std_logic;                      -- sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	signal sdram_s1_translator_avalon_anti_slave_0_byteenable                                           : std_logic_vector(1 downto 0);   -- sdram_s1_translator:av_byteenable -> sdram_s1_translator_avalon_anti_slave_0_byteenable:in
	signal system_id_control_slave_translator_avalon_anti_slave_0_address                               : std_logic_vector(0 downto 0);   -- system_id_control_slave_translator:av_address -> system_id:address
	signal system_id_control_slave_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0);  -- system_id:readdata -> system_id_control_slave_translator:av_readdata
	signal pll_pll_slave_translator_avalon_anti_slave_0_writedata                                       : std_logic_vector(31 downto 0);  -- pll_pll_slave_translator:av_writedata -> pll:writedata
	signal pll_pll_slave_translator_avalon_anti_slave_0_address                                         : std_logic_vector(1 downto 0);   -- pll_pll_slave_translator:av_address -> pll:address
	signal pll_pll_slave_translator_avalon_anti_slave_0_write                                           : std_logic;                      -- pll_pll_slave_translator:av_write -> pll:write
	signal pll_pll_slave_translator_avalon_anti_slave_0_read                                            : std_logic;                      -- pll_pll_slave_translator:av_read -> pll:read
	signal pll_pll_slave_translator_avalon_anti_slave_0_readdata                                        : std_logic_vector(31 downto 0);  -- pll:readdata -> pll_pll_slave_translator:av_readdata
	signal uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                            : std_logic;                      -- uart:av_waitrequest -> uart_avalon_jtag_slave_translator:av_waitrequest
	signal uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                              : std_logic_vector(31 downto 0);  -- uart_avalon_jtag_slave_translator:av_writedata -> uart:av_writedata
	signal uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address                                : std_logic_vector(0 downto 0);   -- uart_avalon_jtag_slave_translator:av_address -> uart:av_address
	signal uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                             : std_logic;                      -- uart_avalon_jtag_slave_translator:av_chipselect -> uart:av_chipselect
	signal uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                  : std_logic;                      -- uart_avalon_jtag_slave_translator:av_write -> uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                   : std_logic;                      -- uart_avalon_jtag_slave_translator:av_read -> uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                               : std_logic_vector(31 downto 0);  -- uart:av_readdata -> uart_avalon_jtag_slave_translator:av_readdata
	signal timer_0_s1_translator_avalon_anti_slave_0_writedata                                          : std_logic_vector(15 downto 0);  -- timer_0_s1_translator:av_writedata -> timer_0:writedata
	signal timer_0_s1_translator_avalon_anti_slave_0_address                                            : std_logic_vector(2 downto 0);   -- timer_0_s1_translator:av_address -> timer_0:address
	signal timer_0_s1_translator_avalon_anti_slave_0_chipselect                                         : std_logic;                      -- timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	signal timer_0_s1_translator_avalon_anti_slave_0_write                                              : std_logic;                      -- timer_0_s1_translator:av_write -> timer_0_s1_translator_avalon_anti_slave_0_write:in
	signal timer_0_s1_translator_avalon_anti_slave_0_readdata                                           : std_logic_vector(15 downto 0);  -- timer_0:readdata -> timer_0_s1_translator:av_readdata
	signal timer_1_s1_translator_avalon_anti_slave_0_writedata                                          : std_logic_vector(15 downto 0);  -- timer_1_s1_translator:av_writedata -> timer_1:writedata
	signal timer_1_s1_translator_avalon_anti_slave_0_address                                            : std_logic_vector(2 downto 0);   -- timer_1_s1_translator:av_address -> timer_1:address
	signal timer_1_s1_translator_avalon_anti_slave_0_chipselect                                         : std_logic;                      -- timer_1_s1_translator:av_chipselect -> timer_1:chipselect
	signal timer_1_s1_translator_avalon_anti_slave_0_write                                              : std_logic;                      -- timer_1_s1_translator:av_write -> timer_1_s1_translator_avalon_anti_slave_0_write:in
	signal timer_1_s1_translator_avalon_anti_slave_0_readdata                                           : std_logic_vector(15 downto 0);  -- timer_1:readdata -> timer_1_s1_translator:av_readdata
	signal pio_in_sw_s1_translator_avalon_anti_slave_0_address                                          : std_logic_vector(1 downto 0);   -- pio_in_sw_s1_translator:av_address -> pio_in_sw:address
	signal pio_in_sw_s1_translator_avalon_anti_slave_0_readdata                                         : std_logic_vector(31 downto 0);  -- pio_in_sw:readdata -> pio_in_sw_s1_translator:av_readdata
	signal pio_in_key_edge_s1_translator_avalon_anti_slave_0_writedata                                  : std_logic_vector(31 downto 0);  -- pio_in_key_edge_s1_translator:av_writedata -> pio_in_key_edge:writedata
	signal pio_in_key_edge_s1_translator_avalon_anti_slave_0_address                                    : std_logic_vector(1 downto 0);   -- pio_in_key_edge_s1_translator:av_address -> pio_in_key_edge:address
	signal pio_in_key_edge_s1_translator_avalon_anti_slave_0_chipselect                                 : std_logic;                      -- pio_in_key_edge_s1_translator:av_chipselect -> pio_in_key_edge:chipselect
	signal pio_in_key_edge_s1_translator_avalon_anti_slave_0_write                                      : std_logic;                      -- pio_in_key_edge_s1_translator:av_write -> pio_in_key_edge_s1_translator_avalon_anti_slave_0_write:in
	signal pio_in_key_edge_s1_translator_avalon_anti_slave_0_readdata                                   : std_logic_vector(31 downto 0);  -- pio_in_key_edge:readdata -> pio_in_key_edge_s1_translator:av_readdata
	signal pio_in_ext_s1_translator_avalon_anti_slave_0_writedata                                       : std_logic_vector(31 downto 0);  -- pio_in_ext_s1_translator:av_writedata -> pio_in_ext:writedata
	signal pio_in_ext_s1_translator_avalon_anti_slave_0_address                                         : std_logic_vector(1 downto 0);   -- pio_in_ext_s1_translator:av_address -> pio_in_ext:address
	signal pio_in_ext_s1_translator_avalon_anti_slave_0_chipselect                                      : std_logic;                      -- pio_in_ext_s1_translator:av_chipselect -> pio_in_ext:chipselect
	signal pio_in_ext_s1_translator_avalon_anti_slave_0_write                                           : std_logic;                      -- pio_in_ext_s1_translator:av_write -> pio_in_ext_s1_translator_avalon_anti_slave_0_write:in
	signal pio_in_ext_s1_translator_avalon_anti_slave_0_readdata                                        : std_logic_vector(31 downto 0);  -- pio_in_ext:readdata -> pio_in_ext_s1_translator:av_readdata
	signal pio_out_red_s1_translator_avalon_anti_slave_0_writedata                                      : std_logic_vector(31 downto 0);  -- pio_out_red_s1_translator:av_writedata -> pio_out_red:writedata
	signal pio_out_red_s1_translator_avalon_anti_slave_0_address                                        : std_logic_vector(2 downto 0);   -- pio_out_red_s1_translator:av_address -> pio_out_red:address
	signal pio_out_red_s1_translator_avalon_anti_slave_0_chipselect                                     : std_logic;                      -- pio_out_red_s1_translator:av_chipselect -> pio_out_red:chipselect
	signal pio_out_red_s1_translator_avalon_anti_slave_0_write                                          : std_logic;                      -- pio_out_red_s1_translator:av_write -> pio_out_red_s1_translator_avalon_anti_slave_0_write:in
	signal pio_out_red_s1_translator_avalon_anti_slave_0_readdata                                       : std_logic_vector(31 downto 0);  -- pio_out_red:readdata -> pio_out_red_s1_translator:av_readdata
	signal pio_out_green_s1_translator_avalon_anti_slave_0_writedata                                    : std_logic_vector(31 downto 0);  -- pio_out_green_s1_translator:av_writedata -> pio_out_green:writedata
	signal pio_out_green_s1_translator_avalon_anti_slave_0_address                                      : std_logic_vector(2 downto 0);   -- pio_out_green_s1_translator:av_address -> pio_out_green:address
	signal pio_out_green_s1_translator_avalon_anti_slave_0_chipselect                                   : std_logic;                      -- pio_out_green_s1_translator:av_chipselect -> pio_out_green:chipselect
	signal pio_out_green_s1_translator_avalon_anti_slave_0_write                                        : std_logic;                      -- pio_out_green_s1_translator:av_write -> pio_out_green_s1_translator_avalon_anti_slave_0_write:in
	signal pio_out_green_s1_translator_avalon_anti_slave_0_readdata                                     : std_logic_vector(31 downto 0);  -- pio_out_green:readdata -> pio_out_green_s1_translator:av_readdata
	signal pio_out_ext_s1_translator_avalon_anti_slave_0_writedata                                      : std_logic_vector(31 downto 0);  -- pio_out_ext_s1_translator:av_writedata -> pio_out_ext:writedata
	signal pio_out_ext_s1_translator_avalon_anti_slave_0_address                                        : std_logic_vector(2 downto 0);   -- pio_out_ext_s1_translator:av_address -> pio_out_ext:address
	signal pio_out_ext_s1_translator_avalon_anti_slave_0_chipselect                                     : std_logic;                      -- pio_out_ext_s1_translator:av_chipselect -> pio_out_ext:chipselect
	signal pio_out_ext_s1_translator_avalon_anti_slave_0_write                                          : std_logic;                      -- pio_out_ext_s1_translator:av_write -> pio_out_ext_s1_translator_avalon_anti_slave_0_write:in
	signal pio_out_ext_s1_translator_avalon_anti_slave_0_readdata                                       : std_logic_vector(31 downto 0);  -- pio_out_ext:readdata -> pio_out_ext_s1_translator:av_readdata
	signal pio_async_reset_s1_translator_avalon_anti_slave_0_writedata                                  : std_logic_vector(31 downto 0);  -- pio_async_reset_s1_translator:av_writedata -> pio_async_reset:writedata
	signal pio_async_reset_s1_translator_avalon_anti_slave_0_address                                    : std_logic_vector(2 downto 0);   -- pio_async_reset_s1_translator:av_address -> pio_async_reset:address
	signal pio_async_reset_s1_translator_avalon_anti_slave_0_chipselect                                 : std_logic;                      -- pio_async_reset_s1_translator:av_chipselect -> pio_async_reset:chipselect
	signal pio_async_reset_s1_translator_avalon_anti_slave_0_write                                      : std_logic;                      -- pio_async_reset_s1_translator:av_write -> pio_async_reset_s1_translator_avalon_anti_slave_0_write:in
	signal pio_async_reset_s1_translator_avalon_anti_slave_0_readdata                                   : std_logic_vector(31 downto 0);  -- pio_async_reset:readdata -> pio_async_reset_s1_translator:av_readdata
	signal pio_en_mux_s1_translator_avalon_anti_slave_0_writedata                                       : std_logic_vector(31 downto 0);  -- pio_en_mux_s1_translator:av_writedata -> pio_en_mux:writedata
	signal pio_en_mux_s1_translator_avalon_anti_slave_0_address                                         : std_logic_vector(2 downto 0);   -- pio_en_mux_s1_translator:av_address -> pio_en_mux:address
	signal pio_en_mux_s1_translator_avalon_anti_slave_0_chipselect                                      : std_logic;                      -- pio_en_mux_s1_translator:av_chipselect -> pio_en_mux:chipselect
	signal pio_en_mux_s1_translator_avalon_anti_slave_0_write                                           : std_logic;                      -- pio_en_mux_s1_translator:av_write -> pio_en_mux_s1_translator_avalon_anti_slave_0_write:in
	signal pio_en_mux_s1_translator_avalon_anti_slave_0_readdata                                        : std_logic_vector(31 downto 0);  -- pio_en_mux:readdata -> pio_en_mux_s1_translator:av_readdata
	signal pio_direc_s1_translator_avalon_anti_slave_0_writedata                                        : std_logic_vector(31 downto 0);  -- pio_direc_s1_translator:av_writedata -> pio_direc:writedata
	signal pio_direc_s1_translator_avalon_anti_slave_0_address                                          : std_logic_vector(2 downto 0);   -- pio_direc_s1_translator:av_address -> pio_direc:address
	signal pio_direc_s1_translator_avalon_anti_slave_0_chipselect                                       : std_logic;                      -- pio_direc_s1_translator:av_chipselect -> pio_direc:chipselect
	signal pio_direc_s1_translator_avalon_anti_slave_0_write                                            : std_logic;                      -- pio_direc_s1_translator:av_write -> pio_direc_s1_translator_avalon_anti_slave_0_write:in
	signal pio_direc_s1_translator_avalon_anti_slave_0_readdata                                         : std_logic_vector(31 downto 0);  -- pio_direc:readdata -> pio_direc_s1_translator:av_readdata
	signal pio_direc_ram_s1_translator_avalon_anti_slave_0_writedata                                    : std_logic_vector(31 downto 0);  -- pio_direc_ram_s1_translator:av_writedata -> pio_direc_ram:writedata
	signal pio_direc_ram_s1_translator_avalon_anti_slave_0_address                                      : std_logic_vector(2 downto 0);   -- pio_direc_ram_s1_translator:av_address -> pio_direc_ram:address
	signal pio_direc_ram_s1_translator_avalon_anti_slave_0_chipselect                                   : std_logic;                      -- pio_direc_ram_s1_translator:av_chipselect -> pio_direc_ram:chipselect
	signal pio_direc_ram_s1_translator_avalon_anti_slave_0_write                                        : std_logic;                      -- pio_direc_ram_s1_translator:av_write -> pio_direc_ram_s1_translator_avalon_anti_slave_0_write:in
	signal pio_direc_ram_s1_translator_avalon_anti_slave_0_readdata                                     : std_logic_vector(31 downto 0);  -- pio_direc_ram:readdata -> pio_direc_ram_s1_translator:av_readdata
	signal pio_wr_s1_translator_avalon_anti_slave_0_writedata                                           : std_logic_vector(31 downto 0);  -- pio_wr_s1_translator:av_writedata -> pio_wr:writedata
	signal pio_wr_s1_translator_avalon_anti_slave_0_address                                             : std_logic_vector(2 downto 0);   -- pio_wr_s1_translator:av_address -> pio_wr:address
	signal pio_wr_s1_translator_avalon_anti_slave_0_chipselect                                          : std_logic;                      -- pio_wr_s1_translator:av_chipselect -> pio_wr:chipselect
	signal pio_wr_s1_translator_avalon_anti_slave_0_write                                               : std_logic;                      -- pio_wr_s1_translator:av_write -> pio_wr_s1_translator_avalon_anti_slave_0_write:in
	signal pio_wr_s1_translator_avalon_anti_slave_0_readdata                                            : std_logic_vector(31 downto 0);  -- pio_wr:readdata -> pio_wr_s1_translator:av_readdata
	signal pio_sel_salida_s1_translator_avalon_anti_slave_0_writedata                                   : std_logic_vector(31 downto 0);  -- pio_sel_salida_s1_translator:av_writedata -> pio_sel_salida:writedata
	signal pio_sel_salida_s1_translator_avalon_anti_slave_0_address                                     : std_logic_vector(2 downto 0);   -- pio_sel_salida_s1_translator:av_address -> pio_sel_salida:address
	signal pio_sel_salida_s1_translator_avalon_anti_slave_0_chipselect                                  : std_logic;                      -- pio_sel_salida_s1_translator:av_chipselect -> pio_sel_salida:chipselect
	signal pio_sel_salida_s1_translator_avalon_anti_slave_0_write                                       : std_logic;                      -- pio_sel_salida_s1_translator:av_write -> pio_sel_salida_s1_translator_avalon_anti_slave_0_write:in
	signal pio_sel_salida_s1_translator_avalon_anti_slave_0_readdata                                    : std_logic_vector(31 downto 0);  -- pio_sel_salida:readdata -> pio_sel_salida_s1_translator:av_readdata
	signal pio_datos_s1_translator_avalon_anti_slave_0_writedata                                        : std_logic_vector(31 downto 0);  -- pio_datos_s1_translator:av_writedata -> pio_datos:writedata
	signal pio_datos_s1_translator_avalon_anti_slave_0_address                                          : std_logic_vector(2 downto 0);   -- pio_datos_s1_translator:av_address -> pio_datos:address
	signal pio_datos_s1_translator_avalon_anti_slave_0_chipselect                                       : std_logic;                      -- pio_datos_s1_translator:av_chipselect -> pio_datos:chipselect
	signal pio_datos_s1_translator_avalon_anti_slave_0_write                                            : std_logic;                      -- pio_datos_s1_translator:av_write -> pio_datos_s1_translator_avalon_anti_slave_0_write:in
	signal pio_datos_s1_translator_avalon_anti_slave_0_readdata                                         : std_logic_vector(31 downto 0);  -- pio_datos:readdata -> pio_datos_s1_translator:av_readdata
	signal pio_compara_int_0_s1_translator_avalon_anti_slave_0_writedata                                : std_logic_vector(31 downto 0);  -- pio_compara_int_0_s1_translator:av_writedata -> pio_compara_int_0:writedata
	signal pio_compara_int_0_s1_translator_avalon_anti_slave_0_address                                  : std_logic_vector(1 downto 0);   -- pio_compara_int_0_s1_translator:av_address -> pio_compara_int_0:address
	signal pio_compara_int_0_s1_translator_avalon_anti_slave_0_chipselect                               : std_logic;                      -- pio_compara_int_0_s1_translator:av_chipselect -> pio_compara_int_0:chipselect
	signal pio_compara_int_0_s1_translator_avalon_anti_slave_0_write                                    : std_logic;                      -- pio_compara_int_0_s1_translator:av_write -> pio_compara_int_0_s1_translator_avalon_anti_slave_0_write:in
	signal pio_compara_int_0_s1_translator_avalon_anti_slave_0_readdata                                 : std_logic_vector(31 downto 0);  -- pio_compara_int_0:readdata -> pio_compara_int_0_s1_translator:av_readdata
	signal pio_compara_int_1_s1_translator_avalon_anti_slave_0_writedata                                : std_logic_vector(31 downto 0);  -- pio_compara_int_1_s1_translator:av_writedata -> pio_compara_int_1:writedata
	signal pio_compara_int_1_s1_translator_avalon_anti_slave_0_address                                  : std_logic_vector(1 downto 0);   -- pio_compara_int_1_s1_translator:av_address -> pio_compara_int_1:address
	signal pio_compara_int_1_s1_translator_avalon_anti_slave_0_chipselect                               : std_logic;                      -- pio_compara_int_1_s1_translator:av_chipselect -> pio_compara_int_1:chipselect
	signal pio_compara_int_1_s1_translator_avalon_anti_slave_0_write                                    : std_logic;                      -- pio_compara_int_1_s1_translator:av_write -> pio_compara_int_1_s1_translator_avalon_anti_slave_0_write:in
	signal pio_compara_int_1_s1_translator_avalon_anti_slave_0_readdata                                 : std_logic_vector(31 downto 0);  -- pio_compara_int_1:readdata -> pio_compara_int_1_s1_translator:av_readdata
	signal pio_compara_int_2_s1_translator_avalon_anti_slave_0_writedata                                : std_logic_vector(31 downto 0);  -- pio_compara_int_2_s1_translator:av_writedata -> pio_compara_int_2:writedata
	signal pio_compara_int_2_s1_translator_avalon_anti_slave_0_address                                  : std_logic_vector(1 downto 0);   -- pio_compara_int_2_s1_translator:av_address -> pio_compara_int_2:address
	signal pio_compara_int_2_s1_translator_avalon_anti_slave_0_chipselect                               : std_logic;                      -- pio_compara_int_2_s1_translator:av_chipselect -> pio_compara_int_2:chipselect
	signal pio_compara_int_2_s1_translator_avalon_anti_slave_0_write                                    : std_logic;                      -- pio_compara_int_2_s1_translator:av_write -> pio_compara_int_2_s1_translator_avalon_anti_slave_0_write:in
	signal pio_compara_int_2_s1_translator_avalon_anti_slave_0_readdata                                 : std_logic_vector(31 downto 0);  -- pio_compara_int_2:readdata -> pio_compara_int_2_s1_translator:av_readdata
	signal pio_compara_int_3_s1_translator_avalon_anti_slave_0_writedata                                : std_logic_vector(31 downto 0);  -- pio_compara_int_3_s1_translator:av_writedata -> pio_compara_int_3:writedata
	signal pio_compara_int_3_s1_translator_avalon_anti_slave_0_address                                  : std_logic_vector(1 downto 0);   -- pio_compara_int_3_s1_translator:av_address -> pio_compara_int_3:address
	signal pio_compara_int_3_s1_translator_avalon_anti_slave_0_chipselect                               : std_logic;                      -- pio_compara_int_3_s1_translator:av_chipselect -> pio_compara_int_3:chipselect
	signal pio_compara_int_3_s1_translator_avalon_anti_slave_0_write                                    : std_logic;                      -- pio_compara_int_3_s1_translator:av_write -> pio_compara_int_3_s1_translator_avalon_anti_slave_0_write:in
	signal pio_compara_int_3_s1_translator_avalon_anti_slave_0_readdata                                 : std_logic_vector(31 downto 0);  -- pio_compara_int_3:readdata -> pio_compara_int_3_s1_translator:av_readdata
	signal pio_compara_int_4_s1_translator_avalon_anti_slave_0_writedata                                : std_logic_vector(31 downto 0);  -- pio_compara_int_4_s1_translator:av_writedata -> pio_compara_int_4:writedata
	signal pio_compara_int_4_s1_translator_avalon_anti_slave_0_address                                  : std_logic_vector(1 downto 0);   -- pio_compara_int_4_s1_translator:av_address -> pio_compara_int_4:address
	signal pio_compara_int_4_s1_translator_avalon_anti_slave_0_chipselect                               : std_logic;                      -- pio_compara_int_4_s1_translator:av_chipselect -> pio_compara_int_4:chipselect
	signal pio_compara_int_4_s1_translator_avalon_anti_slave_0_write                                    : std_logic;                      -- pio_compara_int_4_s1_translator:av_write -> pio_compara_int_4_s1_translator_avalon_anti_slave_0_write:in
	signal pio_compara_int_4_s1_translator_avalon_anti_slave_0_readdata                                 : std_logic_vector(31 downto 0);  -- pio_compara_int_4:readdata -> pio_compara_int_4_s1_translator:av_readdata
	signal pio_captura_0_s1_translator_avalon_anti_slave_0_writedata                                    : std_logic_vector(31 downto 0);  -- pio_captura_0_s1_translator:av_writedata -> pio_captura_0:writedata
	signal pio_captura_0_s1_translator_avalon_anti_slave_0_address                                      : std_logic_vector(1 downto 0);   -- pio_captura_0_s1_translator:av_address -> pio_captura_0:address
	signal pio_captura_0_s1_translator_avalon_anti_slave_0_chipselect                                   : std_logic;                      -- pio_captura_0_s1_translator:av_chipselect -> pio_captura_0:chipselect
	signal pio_captura_0_s1_translator_avalon_anti_slave_0_write                                        : std_logic;                      -- pio_captura_0_s1_translator:av_write -> pio_captura_0_s1_translator_avalon_anti_slave_0_write:in
	signal pio_captura_0_s1_translator_avalon_anti_slave_0_readdata                                     : std_logic_vector(31 downto 0);  -- pio_captura_0:readdata -> pio_captura_0_s1_translator:av_readdata
	signal pio_captura_1_s1_translator_avalon_anti_slave_0_writedata                                    : std_logic_vector(31 downto 0);  -- pio_captura_1_s1_translator:av_writedata -> pio_captura_1:writedata
	signal pio_captura_1_s1_translator_avalon_anti_slave_0_address                                      : std_logic_vector(1 downto 0);   -- pio_captura_1_s1_translator:av_address -> pio_captura_1:address
	signal pio_captura_1_s1_translator_avalon_anti_slave_0_chipselect                                   : std_logic;                      -- pio_captura_1_s1_translator:av_chipselect -> pio_captura_1:chipselect
	signal pio_captura_1_s1_translator_avalon_anti_slave_0_write                                        : std_logic;                      -- pio_captura_1_s1_translator:av_write -> pio_captura_1_s1_translator_avalon_anti_slave_0_write:in
	signal pio_captura_1_s1_translator_avalon_anti_slave_0_readdata                                     : std_logic_vector(31 downto 0);  -- pio_captura_1:readdata -> pio_captura_1_s1_translator:av_readdata
	signal pio_captura_2_s1_translator_avalon_anti_slave_0_writedata                                    : std_logic_vector(31 downto 0);  -- pio_captura_2_s1_translator:av_writedata -> pio_captura_2:writedata
	signal pio_captura_2_s1_translator_avalon_anti_slave_0_address                                      : std_logic_vector(1 downto 0);   -- pio_captura_2_s1_translator:av_address -> pio_captura_2:address
	signal pio_captura_2_s1_translator_avalon_anti_slave_0_chipselect                                   : std_logic;                      -- pio_captura_2_s1_translator:av_chipselect -> pio_captura_2:chipselect
	signal pio_captura_2_s1_translator_avalon_anti_slave_0_write                                        : std_logic;                      -- pio_captura_2_s1_translator:av_write -> pio_captura_2_s1_translator_avalon_anti_slave_0_write:in
	signal pio_captura_2_s1_translator_avalon_anti_slave_0_readdata                                     : std_logic_vector(31 downto 0);  -- pio_captura_2:readdata -> pio_captura_2_s1_translator:av_readdata
	signal pio_captura_3_s1_translator_avalon_anti_slave_0_writedata                                    : std_logic_vector(31 downto 0);  -- pio_captura_3_s1_translator:av_writedata -> pio_captura_3:writedata
	signal pio_captura_3_s1_translator_avalon_anti_slave_0_address                                      : std_logic_vector(1 downto 0);   -- pio_captura_3_s1_translator:av_address -> pio_captura_3:address
	signal pio_captura_3_s1_translator_avalon_anti_slave_0_chipselect                                   : std_logic;                      -- pio_captura_3_s1_translator:av_chipselect -> pio_captura_3:chipselect
	signal pio_captura_3_s1_translator_avalon_anti_slave_0_write                                        : std_logic;                      -- pio_captura_3_s1_translator:av_write -> pio_captura_3_s1_translator_avalon_anti_slave_0_write:in
	signal pio_captura_3_s1_translator_avalon_anti_slave_0_readdata                                     : std_logic_vector(31 downto 0);  -- pio_captura_3:readdata -> pio_captura_3_s1_translator:av_readdata
	signal pio_captura_4_s1_translator_avalon_anti_slave_0_writedata                                    : std_logic_vector(31 downto 0);  -- pio_captura_4_s1_translator:av_writedata -> pio_captura_4:writedata
	signal pio_captura_4_s1_translator_avalon_anti_slave_0_address                                      : std_logic_vector(1 downto 0);   -- pio_captura_4_s1_translator:av_address -> pio_captura_4:address
	signal pio_captura_4_s1_translator_avalon_anti_slave_0_chipselect                                   : std_logic;                      -- pio_captura_4_s1_translator:av_chipselect -> pio_captura_4:chipselect
	signal pio_captura_4_s1_translator_avalon_anti_slave_0_write                                        : std_logic;                      -- pio_captura_4_s1_translator:av_write -> pio_captura_4_s1_translator_avalon_anti_slave_0_write:in
	signal pio_captura_4_s1_translator_avalon_anti_slave_0_readdata                                     : std_logic_vector(31 downto 0);  -- pio_captura_4:readdata -> pio_captura_4_s1_translator:av_readdata
	signal pio_in_32_s1_translator_avalon_anti_slave_0_writedata                                        : std_logic_vector(31 downto 0);  -- pio_in_32_s1_translator:av_writedata -> pio_in_32:writedata
	signal pio_in_32_s1_translator_avalon_anti_slave_0_address                                          : std_logic_vector(1 downto 0);   -- pio_in_32_s1_translator:av_address -> pio_in_32:address
	signal pio_in_32_s1_translator_avalon_anti_slave_0_chipselect                                       : std_logic;                      -- pio_in_32_s1_translator:av_chipselect -> pio_in_32:chipselect
	signal pio_in_32_s1_translator_avalon_anti_slave_0_write                                            : std_logic;                      -- pio_in_32_s1_translator:av_write -> pio_in_32_s1_translator_avalon_anti_slave_0_write:in
	signal pio_in_32_s1_translator_avalon_anti_slave_0_readdata                                         : std_logic_vector(31 downto 0);  -- pio_in_32:readdata -> pio_in_32_s1_translator:av_readdata
	signal lcd_control_slave_translator_avalon_anti_slave_0_writedata                                   : std_logic_vector(7 downto 0);   -- lcd_control_slave_translator:av_writedata -> lcd:writedata
	signal lcd_control_slave_translator_avalon_anti_slave_0_address                                     : std_logic_vector(1 downto 0);   -- lcd_control_slave_translator:av_address -> lcd:address
	signal lcd_control_slave_translator_avalon_anti_slave_0_write                                       : std_logic;                      -- lcd_control_slave_translator:av_write -> lcd:write
	signal lcd_control_slave_translator_avalon_anti_slave_0_read                                        : std_logic;                      -- lcd_control_slave_translator:av_read -> lcd:read
	signal lcd_control_slave_translator_avalon_anti_slave_0_readdata                                    : std_logic_vector(7 downto 0);   -- lcd:readdata -> lcd_control_slave_translator:av_readdata
	signal lcd_control_slave_translator_avalon_anti_slave_0_begintransfer                               : std_logic;                      -- lcd_control_slave_translator:av_begintransfer -> lcd:begintransfer
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_writedata                              : std_logic_vector(15 downto 0);  -- DM9000A_avalon_slave_0_translator:av_writedata -> DM9000A:iDATA
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_address                                : std_logic_vector(0 downto 0);   -- DM9000A_avalon_slave_0_translator:av_address -> DM9000A:iCMD
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect                             : std_logic;                      -- DM9000A_avalon_slave_0_translator:av_chipselect -> dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect:in
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write                                  : std_logic;                      -- DM9000A_avalon_slave_0_translator:av_write -> dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write:in
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read                                   : std_logic;                      -- DM9000A_avalon_slave_0_translator:av_read -> dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read:in
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_readdata                               : std_logic_vector(15 downto 0);  -- DM9000A:oDATA -> DM9000A_avalon_slave_0_translator:av_readdata
	signal cpu_instruction_master_translator_avalon_universal_master_0_waitrequest                      : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_instruction_master_translator:uav_waitrequest
	signal cpu_instruction_master_translator_avalon_universal_master_0_burstcount                       : std_logic_vector(2 downto 0);   -- cpu_instruction_master_translator:uav_burstcount -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_instruction_master_translator_avalon_universal_master_0_writedata                        : std_logic_vector(31 downto 0);  -- cpu_instruction_master_translator:uav_writedata -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_instruction_master_translator_avalon_universal_master_0_address                          : std_logic_vector(24 downto 0);  -- cpu_instruction_master_translator:uav_address -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal cpu_instruction_master_translator_avalon_universal_master_0_lock                             : std_logic;                      -- cpu_instruction_master_translator:uav_lock -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_instruction_master_translator_avalon_universal_master_0_write                            : std_logic;                      -- cpu_instruction_master_translator:uav_write -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal cpu_instruction_master_translator_avalon_universal_master_0_read                             : std_logic;                      -- cpu_instruction_master_translator:uav_read -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal cpu_instruction_master_translator_avalon_universal_master_0_readdata                         : std_logic_vector(31 downto 0);  -- cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_instruction_master_translator:uav_readdata
	signal cpu_instruction_master_translator_avalon_universal_master_0_debugaccess                      : std_logic;                      -- cpu_instruction_master_translator:uav_debugaccess -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_instruction_master_translator_avalon_universal_master_0_byteenable                       : std_logic_vector(3 downto 0);   -- cpu_instruction_master_translator:uav_byteenable -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid                    : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_instruction_master_translator:uav_readdatavalid
	signal cpu_data_master_translator_avalon_universal_master_0_waitrequest                             : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_data_master_translator:uav_waitrequest
	signal cpu_data_master_translator_avalon_universal_master_0_burstcount                              : std_logic_vector(2 downto 0);   -- cpu_data_master_translator:uav_burstcount -> cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_data_master_translator_avalon_universal_master_0_writedata                               : std_logic_vector(31 downto 0);  -- cpu_data_master_translator:uav_writedata -> cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_data_master_translator_avalon_universal_master_0_address                                 : std_logic_vector(24 downto 0);  -- cpu_data_master_translator:uav_address -> cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	signal cpu_data_master_translator_avalon_universal_master_0_lock                                    : std_logic;                      -- cpu_data_master_translator:uav_lock -> cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_data_master_translator_avalon_universal_master_0_write                                   : std_logic;                      -- cpu_data_master_translator:uav_write -> cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	signal cpu_data_master_translator_avalon_universal_master_0_read                                    : std_logic;                      -- cpu_data_master_translator:uav_read -> cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	signal cpu_data_master_translator_avalon_universal_master_0_readdata                                : std_logic_vector(31 downto 0);  -- cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_data_master_translator:uav_readdata
	signal cpu_data_master_translator_avalon_universal_master_0_debugaccess                             : std_logic;                      -- cpu_data_master_translator:uav_debugaccess -> cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_data_master_translator_avalon_universal_master_0_byteenable                              : std_logic_vector(3 downto 0);   -- cpu_data_master_translator:uav_byteenable -> cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_data_master_translator_avalon_universal_master_0_readdatavalid                           : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_data_master_translator:uav_readdatavalid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest               : std_logic;                      -- cpu_jtag_debug_module_translator:uav_waitrequest -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount                : std_logic_vector(2 downto 0);   -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_jtag_debug_module_translator:uav_burstcount
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata                 : std_logic_vector(31 downto 0);  -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_jtag_debug_module_translator:uav_writedata
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                   : std_logic_vector(24 downto 0);  -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_jtag_debug_module_translator:uav_address
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                     : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_jtag_debug_module_translator:uav_write
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                      : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_jtag_debug_module_translator:uav_lock
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                      : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_jtag_debug_module_translator:uav_read
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                  : std_logic_vector(31 downto 0);  -- cpu_jtag_debug_module_translator:uav_readdata -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid             : std_logic;                      -- cpu_jtag_debug_module_translator:uav_readdatavalid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess               : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_jtag_debug_module_translator:uav_debugaccess
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable                : std_logic_vector(3 downto 0);   -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_jtag_debug_module_translator:uav_byteenable
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket        : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid              : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket      : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data               : std_logic_vector(104 downto 0); -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready              : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket     : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid           : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket   : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data            : std_logic_vector(104 downto 0); -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready           : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid         : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data          : std_logic_vector(33 downto 0);  -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready         : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                            : std_logic;                      -- sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                             : std_logic_vector(1 downto 0);   -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata                              : std_logic_vector(15 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_address                                : std_logic_vector(24 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_write                                  : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock                                   : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_read                                   : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata                               : std_logic_vector(15 downto 0);  -- sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                          : std_logic;                      -- sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                            : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	signal sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                             : std_logic_vector(1 downto 0);   -- sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                     : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                           : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                   : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data                            : std_logic_vector(86 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                           : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                  : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                        : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                         : std_logic_vector(86 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                        : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                      : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                       : std_logic_vector(17 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                      : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                      : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                       : std_logic_vector(17 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                      : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                      -- system_id_control_slave_translator:uav_waitrequest -> system_id_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);   -- system_id_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> system_id_control_slave_translator:uav_burstcount
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0);  -- system_id_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> system_id_control_slave_translator:uav_writedata
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(24 downto 0);  -- system_id_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> system_id_control_slave_translator:uav_address
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> system_id_control_slave_translator:uav_write
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> system_id_control_slave_translator:uav_lock
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> system_id_control_slave_translator:uav_read
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0);  -- system_id_control_slave_translator:uav_readdata -> system_id_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                      -- system_id_control_slave_translator:uav_readdatavalid -> system_id_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> system_id_control_slave_translator:uav_debugaccess
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);   -- system_id_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> system_id_control_slave_translator:uav_byteenable
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(104 downto 0); -- system_id_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> system_id_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> system_id_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> system_id_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> system_id_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(104 downto 0); -- system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> system_id_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> system_id_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0);  -- system_id_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> system_id_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> system_id_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                       : std_logic;                      -- pll_pll_slave_translator:uav_waitrequest -> pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                        : std_logic_vector(2 downto 0);   -- pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> pll_pll_slave_translator:uav_burstcount
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata                         : std_logic_vector(31 downto 0);  -- pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> pll_pll_slave_translator:uav_writedata
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address                           : std_logic_vector(24 downto 0);  -- pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> pll_pll_slave_translator:uav_address
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write                             : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> pll_pll_slave_translator:uav_write
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock                              : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> pll_pll_slave_translator:uav_lock
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read                              : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> pll_pll_slave_translator:uav_read
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata                          : std_logic_vector(31 downto 0);  -- pll_pll_slave_translator:uav_readdata -> pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                     : std_logic;                      -- pll_pll_slave_translator:uav_readdatavalid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                       : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pll_pll_slave_translator:uav_debugaccess
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                        : std_logic_vector(3 downto 0);   -- pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> pll_pll_slave_translator:uav_byteenable
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                      : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket              : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data                       : std_logic_vector(104 downto 0); -- pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                      : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket             : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                   : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket           : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                    : std_logic_vector(104 downto 0); -- pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                   : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                 : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                  : std_logic_vector(33 downto 0);  -- pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                 : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                 : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                  : std_logic_vector(33 downto 0);  -- pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                 : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest              : std_logic;                      -- uart_avalon_jtag_slave_translator:uav_waitrequest -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount               : std_logic_vector(2 downto 0);   -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart_avalon_jtag_slave_translator:uav_burstcount
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata                : std_logic_vector(31 downto 0);  -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> uart_avalon_jtag_slave_translator:uav_writedata
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                  : std_logic_vector(24 downto 0);  -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> uart_avalon_jtag_slave_translator:uav_address
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                    : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> uart_avalon_jtag_slave_translator:uav_write
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                     : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> uart_avalon_jtag_slave_translator:uav_lock
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                     : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> uart_avalon_jtag_slave_translator:uav_read
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                 : std_logic_vector(31 downto 0);  -- uart_avalon_jtag_slave_translator:uav_readdata -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid            : std_logic;                      -- uart_avalon_jtag_slave_translator:uav_readdatavalid -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess              : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart_avalon_jtag_slave_translator:uav_debugaccess
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable               : std_logic_vector(3 downto 0);   -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart_avalon_jtag_slave_translator:uav_byteenable
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket       : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid             : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket     : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data              : std_logic_vector(104 downto 0); -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready             : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid          : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket  : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data           : std_logic_vector(104 downto 0); -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready          : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid        : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         : std_logic_vector(33 downto 0);  -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready        : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                          : std_logic;                      -- timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                           : std_logic_vector(2 downto 0);   -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                            : std_logic_vector(31 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address                              : std_logic_vector(24 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write                                : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                                 : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read                                 : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                             : std_logic_vector(31 downto 0);  -- timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                        : std_logic;                      -- timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                          : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                           : std_logic_vector(3 downto 0);   -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                   : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                         : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                 : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                          : std_logic_vector(104 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                         : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                      : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket              : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                       : std_logic_vector(104 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                      : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                    : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                     : std_logic_vector(33 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                    : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                          : std_logic;                      -- timer_1_s1_translator:uav_waitrequest -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                           : std_logic_vector(2 downto 0);   -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_1_s1_translator:uav_burstcount
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata                            : std_logic_vector(31 downto 0);  -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_1_s1_translator:uav_writedata
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address                              : std_logic_vector(24 downto 0);  -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_1_s1_translator:uav_address
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write                                : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_1_s1_translator:uav_write
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock                                 : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_1_s1_translator:uav_lock
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read                                 : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_1_s1_translator:uav_read
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata                             : std_logic_vector(31 downto 0);  -- timer_1_s1_translator:uav_readdata -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                        : std_logic;                      -- timer_1_s1_translator:uav_readdatavalid -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                          : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_1_s1_translator:uav_debugaccess
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                           : std_logic_vector(3 downto 0);   -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_1_s1_translator:uav_byteenable
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                   : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                         : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                 : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data                          : std_logic_vector(104 downto 0); -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                         : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                      : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket              : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                       : std_logic_vector(104 downto 0); -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                      : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                    : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                     : std_logic_vector(33 downto 0);  -- timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                    : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                        : std_logic;                      -- pio_in_sw_s1_translator:uav_waitrequest -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                         : std_logic_vector(2 downto 0);   -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_in_sw_s1_translator:uav_burstcount
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata                          : std_logic_vector(31 downto 0);  -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_in_sw_s1_translator:uav_writedata
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_address                            : std_logic_vector(24 downto 0);  -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_in_sw_s1_translator:uav_address
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_write                              : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_in_sw_s1_translator:uav_write
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_lock                               : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_in_sw_s1_translator:uav_lock
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_read                               : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_in_sw_s1_translator:uav_read
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata                           : std_logic_vector(31 downto 0);  -- pio_in_sw_s1_translator:uav_readdata -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                      : std_logic;                      -- pio_in_sw_s1_translator:uav_readdatavalid -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                        : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_in_sw_s1_translator:uav_debugaccess
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                         : std_logic_vector(3 downto 0);   -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_in_sw_s1_translator:uav_byteenable
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                 : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                       : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket               : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data                        : std_logic_vector(104 downto 0); -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                       : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket              : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                    : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket            : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                     : std_logic_vector(104 downto 0); -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                    : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                  : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                   : std_logic_vector(33 downto 0);  -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                  : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                  : std_logic;                      -- pio_in_key_edge_s1_translator:uav_waitrequest -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                   : std_logic_vector(2 downto 0);   -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_in_key_edge_s1_translator:uav_burstcount
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_writedata                    : std_logic_vector(31 downto 0);  -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_in_key_edge_s1_translator:uav_writedata
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_address                      : std_logic_vector(24 downto 0);  -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_in_key_edge_s1_translator:uav_address
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_write                        : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_in_key_edge_s1_translator:uav_write
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_lock                         : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_in_key_edge_s1_translator:uav_lock
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_read                         : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_in_key_edge_s1_translator:uav_read
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_readdata                     : std_logic_vector(31 downto 0);  -- pio_in_key_edge_s1_translator:uav_readdata -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                : std_logic;                      -- pio_in_key_edge_s1_translator:uav_readdatavalid -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                  : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_in_key_edge_s1_translator:uav_debugaccess
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                   : std_logic_vector(3 downto 0);   -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_in_key_edge_s1_translator:uav_byteenable
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket           : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                 : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket         : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rf_source_data                  : std_logic_vector(104 downto 0); -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                 : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket        : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid              : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket      : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data               : std_logic_vector(104 downto 0); -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready              : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid            : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data             : std_logic_vector(33 downto 0);  -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready            : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                       : std_logic;                      -- pio_in_ext_s1_translator:uav_waitrequest -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                        : std_logic_vector(2 downto 0);   -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_in_ext_s1_translator:uav_burstcount
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_writedata                         : std_logic_vector(31 downto 0);  -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_in_ext_s1_translator:uav_writedata
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_address                           : std_logic_vector(24 downto 0);  -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_in_ext_s1_translator:uav_address
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_write                             : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_in_ext_s1_translator:uav_write
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_lock                              : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_in_ext_s1_translator:uav_lock
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_read                              : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_in_ext_s1_translator:uav_read
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_readdata                          : std_logic_vector(31 downto 0);  -- pio_in_ext_s1_translator:uav_readdata -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                     : std_logic;                      -- pio_in_ext_s1_translator:uav_readdatavalid -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                       : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_in_ext_s1_translator:uav_debugaccess
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                        : std_logic_vector(3 downto 0);   -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_in_ext_s1_translator:uav_byteenable
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                      : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket              : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_data                       : std_logic_vector(104 downto 0); -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                      : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket             : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                   : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket           : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                    : std_logic_vector(104 downto 0); -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                   : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                 : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                  : std_logic_vector(33 downto 0);  -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                 : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                      : std_logic;                      -- pio_out_red_s1_translator:uav_waitrequest -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                       : std_logic_vector(2 downto 0);   -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_out_red_s1_translator:uav_burstcount
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_writedata                        : std_logic_vector(31 downto 0);  -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_out_red_s1_translator:uav_writedata
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_address                          : std_logic_vector(24 downto 0);  -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_out_red_s1_translator:uav_address
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_write                            : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_out_red_s1_translator:uav_write
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_lock                             : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_out_red_s1_translator:uav_lock
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_read                             : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_out_red_s1_translator:uav_read
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_readdata                         : std_logic_vector(31 downto 0);  -- pio_out_red_s1_translator:uav_readdata -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                    : std_logic;                      -- pio_out_red_s1_translator:uav_readdatavalid -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                      : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_out_red_s1_translator:uav_debugaccess
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                       : std_logic_vector(3 downto 0);   -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_out_red_s1_translator:uav_byteenable
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket               : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                     : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket             : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rf_source_data                      : std_logic_vector(104 downto 0); -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                     : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket            : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                  : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket          : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                   : std_logic_vector(104 downto 0); -- pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                  : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                 : std_logic_vector(33 downto 0);  -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                    : std_logic;                      -- pio_out_green_s1_translator:uav_waitrequest -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                     : std_logic_vector(2 downto 0);   -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_out_green_s1_translator:uav_burstcount
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_writedata                      : std_logic_vector(31 downto 0);  -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_out_green_s1_translator:uav_writedata
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_address                        : std_logic_vector(24 downto 0);  -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_out_green_s1_translator:uav_address
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_write                          : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_out_green_s1_translator:uav_write
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_lock                           : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_out_green_s1_translator:uav_lock
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_read                           : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_out_green_s1_translator:uav_read
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_readdata                       : std_logic_vector(31 downto 0);  -- pio_out_green_s1_translator:uav_readdata -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                  : std_logic;                      -- pio_out_green_s1_translator:uav_readdatavalid -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                    : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_out_green_s1_translator:uav_debugaccess
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                     : std_logic_vector(3 downto 0);   -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_out_green_s1_translator:uav_byteenable
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket             : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                   : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket           : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rf_source_data                    : std_logic_vector(104 downto 0); -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                   : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket          : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket        : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                 : std_logic_vector(104 downto 0); -- pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid              : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data               : std_logic_vector(33 downto 0);  -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready              : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                      : std_logic;                      -- pio_out_ext_s1_translator:uav_waitrequest -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                       : std_logic_vector(2 downto 0);   -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_out_ext_s1_translator:uav_burstcount
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_writedata                        : std_logic_vector(31 downto 0);  -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_out_ext_s1_translator:uav_writedata
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_address                          : std_logic_vector(24 downto 0);  -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_out_ext_s1_translator:uav_address
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_write                            : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_out_ext_s1_translator:uav_write
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_lock                             : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_out_ext_s1_translator:uav_lock
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_read                             : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_out_ext_s1_translator:uav_read
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_readdata                         : std_logic_vector(31 downto 0);  -- pio_out_ext_s1_translator:uav_readdata -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                    : std_logic;                      -- pio_out_ext_s1_translator:uav_readdatavalid -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                      : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_out_ext_s1_translator:uav_debugaccess
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                       : std_logic_vector(3 downto 0);   -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_out_ext_s1_translator:uav_byteenable
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket               : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                     : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket             : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_data                      : std_logic_vector(104 downto 0); -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                     : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket            : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                  : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket          : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                   : std_logic_vector(104 downto 0); -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                  : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                 : std_logic_vector(33 downto 0);  -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                  : std_logic;                      -- pio_async_reset_s1_translator:uav_waitrequest -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                   : std_logic_vector(2 downto 0);   -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_async_reset_s1_translator:uav_burstcount
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_writedata                    : std_logic_vector(31 downto 0);  -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_async_reset_s1_translator:uav_writedata
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_address                      : std_logic_vector(24 downto 0);  -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_async_reset_s1_translator:uav_address
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_write                        : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_async_reset_s1_translator:uav_write
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_lock                         : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_async_reset_s1_translator:uav_lock
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_read                         : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_async_reset_s1_translator:uav_read
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_readdata                     : std_logic_vector(31 downto 0);  -- pio_async_reset_s1_translator:uav_readdata -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                : std_logic;                      -- pio_async_reset_s1_translator:uav_readdatavalid -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                  : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_async_reset_s1_translator:uav_debugaccess
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                   : std_logic_vector(3 downto 0);   -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_async_reset_s1_translator:uav_byteenable
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket           : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                 : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket         : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rf_source_data                  : std_logic_vector(104 downto 0); -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                 : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket        : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid              : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket      : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data               : std_logic_vector(104 downto 0); -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready              : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid            : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data             : std_logic_vector(33 downto 0);  -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready            : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                       : std_logic;                      -- pio_en_mux_s1_translator:uav_waitrequest -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                        : std_logic_vector(2 downto 0);   -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_en_mux_s1_translator:uav_burstcount
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_writedata                         : std_logic_vector(31 downto 0);  -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_en_mux_s1_translator:uav_writedata
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_address                           : std_logic_vector(24 downto 0);  -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_en_mux_s1_translator:uav_address
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_write                             : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_en_mux_s1_translator:uav_write
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_lock                              : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_en_mux_s1_translator:uav_lock
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_read                              : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_en_mux_s1_translator:uav_read
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_readdata                          : std_logic_vector(31 downto 0);  -- pio_en_mux_s1_translator:uav_readdata -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                     : std_logic;                      -- pio_en_mux_s1_translator:uav_readdatavalid -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                       : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_en_mux_s1_translator:uav_debugaccess
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                        : std_logic_vector(3 downto 0);   -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_en_mux_s1_translator:uav_byteenable
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                      : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket              : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rf_source_data                       : std_logic_vector(104 downto 0); -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                      : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket             : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                   : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket           : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                    : std_logic_vector(104 downto 0); -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                   : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                 : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                  : std_logic_vector(33 downto 0);  -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                 : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                        : std_logic;                      -- pio_direc_s1_translator:uav_waitrequest -> pio_direc_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                         : std_logic_vector(2 downto 0);   -- pio_direc_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_direc_s1_translator:uav_burstcount
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_writedata                          : std_logic_vector(31 downto 0);  -- pio_direc_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_direc_s1_translator:uav_writedata
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_address                            : std_logic_vector(24 downto 0);  -- pio_direc_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_direc_s1_translator:uav_address
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_write                              : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_direc_s1_translator:uav_write
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_lock                               : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_direc_s1_translator:uav_lock
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_read                               : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_direc_s1_translator:uav_read
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_readdata                           : std_logic_vector(31 downto 0);  -- pio_direc_s1_translator:uav_readdata -> pio_direc_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                      : std_logic;                      -- pio_direc_s1_translator:uav_readdatavalid -> pio_direc_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                        : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_direc_s1_translator:uav_debugaccess
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                         : std_logic_vector(3 downto 0);   -- pio_direc_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_direc_s1_translator:uav_byteenable
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                 : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                       : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket               : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rf_source_data                        : std_logic_vector(104 downto 0); -- pio_direc_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                       : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_direc_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket              : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_direc_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                    : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_direc_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket            : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_direc_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                     : std_logic_vector(104 downto 0); -- pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_direc_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                    : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                  : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_direc_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                   : std_logic_vector(33 downto 0);  -- pio_direc_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_direc_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                  : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_direc_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                    : std_logic;                      -- pio_direc_ram_s1_translator:uav_waitrequest -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                     : std_logic_vector(2 downto 0);   -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_direc_ram_s1_translator:uav_burstcount
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata                      : std_logic_vector(31 downto 0);  -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_direc_ram_s1_translator:uav_writedata
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_address                        : std_logic_vector(24 downto 0);  -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_direc_ram_s1_translator:uav_address
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_write                          : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_direc_ram_s1_translator:uav_write
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock                           : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_direc_ram_s1_translator:uav_lock
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_read                           : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_direc_ram_s1_translator:uav_read
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata                       : std_logic_vector(31 downto 0);  -- pio_direc_ram_s1_translator:uav_readdata -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                  : std_logic;                      -- pio_direc_ram_s1_translator:uav_readdatavalid -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                    : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_direc_ram_s1_translator:uav_debugaccess
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                     : std_logic_vector(3 downto 0);   -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_direc_ram_s1_translator:uav_byteenable
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket             : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                   : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket           : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data                    : std_logic_vector(104 downto 0); -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                   : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket          : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket        : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                 : std_logic_vector(104 downto 0); -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid              : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data               : std_logic_vector(33 downto 0);  -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready              : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                           : std_logic;                      -- pio_wr_s1_translator:uav_waitrequest -> pio_wr_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                            : std_logic_vector(2 downto 0);   -- pio_wr_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_wr_s1_translator:uav_burstcount
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_writedata                             : std_logic_vector(31 downto 0);  -- pio_wr_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_wr_s1_translator:uav_writedata
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_address                               : std_logic_vector(24 downto 0);  -- pio_wr_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_wr_s1_translator:uav_address
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_write                                 : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_wr_s1_translator:uav_write
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_lock                                  : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_wr_s1_translator:uav_lock
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_read                                  : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_wr_s1_translator:uav_read
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_readdata                              : std_logic_vector(31 downto 0);  -- pio_wr_s1_translator:uav_readdata -> pio_wr_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                         : std_logic;                      -- pio_wr_s1_translator:uav_readdatavalid -> pio_wr_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                           : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_wr_s1_translator:uav_debugaccess
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                            : std_logic_vector(3 downto 0);   -- pio_wr_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_wr_s1_translator:uav_byteenable
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                    : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                          : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                  : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rf_source_data                           : std_logic_vector(104 downto 0); -- pio_wr_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                          : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_wr_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                 : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_wr_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                       : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_wr_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket               : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_wr_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                        : std_logic_vector(104 downto 0); -- pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_wr_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                       : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                     : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_wr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                      : std_logic_vector(33 downto 0);  -- pio_wr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_wr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                     : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_wr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                   : std_logic;                      -- pio_sel_salida_s1_translator:uav_waitrequest -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                    : std_logic_vector(2 downto 0);   -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_sel_salida_s1_translator:uav_burstcount
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_writedata                     : std_logic_vector(31 downto 0);  -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_sel_salida_s1_translator:uav_writedata
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_address                       : std_logic_vector(24 downto 0);  -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_sel_salida_s1_translator:uav_address
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_write                         : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_sel_salida_s1_translator:uav_write
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_lock                          : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_sel_salida_s1_translator:uav_lock
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_read                          : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_sel_salida_s1_translator:uav_read
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_readdata                      : std_logic_vector(31 downto 0);  -- pio_sel_salida_s1_translator:uav_readdata -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                 : std_logic;                      -- pio_sel_salida_s1_translator:uav_readdatavalid -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                   : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_sel_salida_s1_translator:uav_debugaccess
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                    : std_logic_vector(3 downto 0);   -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_sel_salida_s1_translator:uav_byteenable
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket            : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                  : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket          : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rf_source_data                   : std_logic_vector(104 downto 0); -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                  : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket         : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid               : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket       : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                : std_logic_vector(104 downto 0); -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready               : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid             : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data              : std_logic_vector(33 downto 0);  -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready             : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                        : std_logic;                      -- pio_datos_s1_translator:uav_waitrequest -> pio_datos_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                         : std_logic_vector(2 downto 0);   -- pio_datos_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_datos_s1_translator:uav_burstcount
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_writedata                          : std_logic_vector(31 downto 0);  -- pio_datos_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_datos_s1_translator:uav_writedata
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_address                            : std_logic_vector(24 downto 0);  -- pio_datos_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_datos_s1_translator:uav_address
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_write                              : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_datos_s1_translator:uav_write
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_lock                               : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_datos_s1_translator:uav_lock
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_read                               : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_datos_s1_translator:uav_read
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_readdata                           : std_logic_vector(31 downto 0);  -- pio_datos_s1_translator:uav_readdata -> pio_datos_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                      : std_logic;                      -- pio_datos_s1_translator:uav_readdatavalid -> pio_datos_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                        : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_datos_s1_translator:uav_debugaccess
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                         : std_logic_vector(3 downto 0);   -- pio_datos_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_datos_s1_translator:uav_byteenable
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                 : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                       : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket               : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rf_source_data                        : std_logic_vector(104 downto 0); -- pio_datos_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                       : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_datos_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket              : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_datos_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                    : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_datos_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket            : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_datos_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                     : std_logic_vector(104 downto 0); -- pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_datos_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                    : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                  : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_datos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                   : std_logic_vector(33 downto 0);  -- pio_datos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_datos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                  : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_datos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                : std_logic;                      -- pio_compara_int_0_s1_translator:uav_waitrequest -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                 : std_logic_vector(2 downto 0);   -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_compara_int_0_s1_translator:uav_burstcount
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                  : std_logic_vector(31 downto 0);  -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_compara_int_0_s1_translator:uav_writedata
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_address                    : std_logic_vector(24 downto 0);  -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_compara_int_0_s1_translator:uav_address
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_write                      : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_compara_int_0_s1_translator:uav_write
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                       : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_compara_int_0_s1_translator:uav_lock
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_read                       : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_compara_int_0_s1_translator:uav_read
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                   : std_logic_vector(31 downto 0);  -- pio_compara_int_0_s1_translator:uav_readdata -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid              : std_logic;                      -- pio_compara_int_0_s1_translator:uav_readdatavalid -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_compara_int_0_s1_translator:uav_debugaccess
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                 : std_logic_vector(3 downto 0);   -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_compara_int_0_s1_translator:uav_byteenable
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket         : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid               : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket       : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                : std_logic_vector(104 downto 0); -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready               : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket      : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid            : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket    : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data             : std_logic_vector(104 downto 0); -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready            : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid          : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data           : std_logic_vector(33 downto 0);  -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready          : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                : std_logic;                      -- pio_compara_int_1_s1_translator:uav_waitrequest -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                 : std_logic_vector(2 downto 0);   -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_compara_int_1_s1_translator:uav_burstcount
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata                  : std_logic_vector(31 downto 0);  -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_compara_int_1_s1_translator:uav_writedata
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_address                    : std_logic_vector(24 downto 0);  -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_compara_int_1_s1_translator:uav_address
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_write                      : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_compara_int_1_s1_translator:uav_write
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_lock                       : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_compara_int_1_s1_translator:uav_lock
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_read                       : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_compara_int_1_s1_translator:uav_read
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata                   : std_logic_vector(31 downto 0);  -- pio_compara_int_1_s1_translator:uav_readdata -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid              : std_logic;                      -- pio_compara_int_1_s1_translator:uav_readdatavalid -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_compara_int_1_s1_translator:uav_debugaccess
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                 : std_logic_vector(3 downto 0);   -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_compara_int_1_s1_translator:uav_byteenable
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket         : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid               : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket       : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data                : std_logic_vector(104 downto 0); -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready               : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket      : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid            : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket    : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data             : std_logic_vector(104 downto 0); -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready            : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid          : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data           : std_logic_vector(33 downto 0);  -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready          : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                : std_logic;                      -- pio_compara_int_2_s1_translator:uav_waitrequest -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                 : std_logic_vector(2 downto 0);   -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_compara_int_2_s1_translator:uav_burstcount
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata                  : std_logic_vector(31 downto 0);  -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_compara_int_2_s1_translator:uav_writedata
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_address                    : std_logic_vector(24 downto 0);  -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_compara_int_2_s1_translator:uav_address
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_write                      : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_compara_int_2_s1_translator:uav_write
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_lock                       : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_compara_int_2_s1_translator:uav_lock
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_read                       : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_compara_int_2_s1_translator:uav_read
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata                   : std_logic_vector(31 downto 0);  -- pio_compara_int_2_s1_translator:uav_readdata -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid              : std_logic;                      -- pio_compara_int_2_s1_translator:uav_readdatavalid -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_compara_int_2_s1_translator:uav_debugaccess
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                 : std_logic_vector(3 downto 0);   -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_compara_int_2_s1_translator:uav_byteenable
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket         : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid               : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket       : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data                : std_logic_vector(104 downto 0); -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready               : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket      : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid            : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket    : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data             : std_logic_vector(104 downto 0); -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready            : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid          : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data           : std_logic_vector(33 downto 0);  -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready          : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                : std_logic;                      -- pio_compara_int_3_s1_translator:uav_waitrequest -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                 : std_logic_vector(2 downto 0);   -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_compara_int_3_s1_translator:uav_burstcount
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata                  : std_logic_vector(31 downto 0);  -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_compara_int_3_s1_translator:uav_writedata
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_address                    : std_logic_vector(24 downto 0);  -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_compara_int_3_s1_translator:uav_address
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_write                      : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_compara_int_3_s1_translator:uav_write
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_lock                       : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_compara_int_3_s1_translator:uav_lock
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_read                       : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_compara_int_3_s1_translator:uav_read
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata                   : std_logic_vector(31 downto 0);  -- pio_compara_int_3_s1_translator:uav_readdata -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid              : std_logic;                      -- pio_compara_int_3_s1_translator:uav_readdatavalid -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_compara_int_3_s1_translator:uav_debugaccess
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                 : std_logic_vector(3 downto 0);   -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_compara_int_3_s1_translator:uav_byteenable
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket         : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid               : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket       : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data                : std_logic_vector(104 downto 0); -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready               : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket      : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid            : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket    : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data             : std_logic_vector(104 downto 0); -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready            : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid          : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data           : std_logic_vector(33 downto 0);  -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready          : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                : std_logic;                      -- pio_compara_int_4_s1_translator:uav_waitrequest -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                 : std_logic_vector(2 downto 0);   -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_compara_int_4_s1_translator:uav_burstcount
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata                  : std_logic_vector(31 downto 0);  -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_compara_int_4_s1_translator:uav_writedata
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_address                    : std_logic_vector(24 downto 0);  -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_compara_int_4_s1_translator:uav_address
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_write                      : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_compara_int_4_s1_translator:uav_write
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_lock                       : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_compara_int_4_s1_translator:uav_lock
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_read                       : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_compara_int_4_s1_translator:uav_read
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata                   : std_logic_vector(31 downto 0);  -- pio_compara_int_4_s1_translator:uav_readdata -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid              : std_logic;                      -- pio_compara_int_4_s1_translator:uav_readdatavalid -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_compara_int_4_s1_translator:uav_debugaccess
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                 : std_logic_vector(3 downto 0);   -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_compara_int_4_s1_translator:uav_byteenable
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket         : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid               : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket       : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data                : std_logic_vector(104 downto 0); -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready               : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket      : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid            : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket    : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data             : std_logic_vector(104 downto 0); -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready            : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid          : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data           : std_logic_vector(33 downto 0);  -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready          : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                    : std_logic;                      -- pio_captura_0_s1_translator:uav_waitrequest -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                     : std_logic_vector(2 downto 0);   -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_captura_0_s1_translator:uav_burstcount
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                      : std_logic_vector(31 downto 0);  -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_captura_0_s1_translator:uav_writedata
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_address                        : std_logic_vector(24 downto 0);  -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_captura_0_s1_translator:uav_address
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_write                          : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_captura_0_s1_translator:uav_write
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                           : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_captura_0_s1_translator:uav_lock
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_read                           : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_captura_0_s1_translator:uav_read
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                       : std_logic_vector(31 downto 0);  -- pio_captura_0_s1_translator:uav_readdata -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                  : std_logic;                      -- pio_captura_0_s1_translator:uav_readdatavalid -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                    : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_captura_0_s1_translator:uav_debugaccess
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                     : std_logic_vector(3 downto 0);   -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_captura_0_s1_translator:uav_byteenable
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket             : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                   : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket           : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                    : std_logic_vector(104 downto 0); -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                   : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket          : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket        : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                 : std_logic_vector(104 downto 0); -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid              : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data               : std_logic_vector(33 downto 0);  -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready              : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                    : std_logic;                      -- pio_captura_1_s1_translator:uav_waitrequest -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                     : std_logic_vector(2 downto 0);   -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_captura_1_s1_translator:uav_burstcount
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata                      : std_logic_vector(31 downto 0);  -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_captura_1_s1_translator:uav_writedata
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_address                        : std_logic_vector(24 downto 0);  -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_captura_1_s1_translator:uav_address
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_write                          : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_captura_1_s1_translator:uav_write
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_lock                           : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_captura_1_s1_translator:uav_lock
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_read                           : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_captura_1_s1_translator:uav_read
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata                       : std_logic_vector(31 downto 0);  -- pio_captura_1_s1_translator:uav_readdata -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                  : std_logic;                      -- pio_captura_1_s1_translator:uav_readdatavalid -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                    : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_captura_1_s1_translator:uav_debugaccess
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                     : std_logic_vector(3 downto 0);   -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_captura_1_s1_translator:uav_byteenable
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket             : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                   : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket           : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data                    : std_logic_vector(104 downto 0); -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                   : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket          : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket        : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                 : std_logic_vector(104 downto 0); -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid              : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data               : std_logic_vector(33 downto 0);  -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready              : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                    : std_logic;                      -- pio_captura_2_s1_translator:uav_waitrequest -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                     : std_logic_vector(2 downto 0);   -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_captura_2_s1_translator:uav_burstcount
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata                      : std_logic_vector(31 downto 0);  -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_captura_2_s1_translator:uav_writedata
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_address                        : std_logic_vector(24 downto 0);  -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_captura_2_s1_translator:uav_address
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_write                          : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_captura_2_s1_translator:uav_write
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_lock                           : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_captura_2_s1_translator:uav_lock
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_read                           : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_captura_2_s1_translator:uav_read
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata                       : std_logic_vector(31 downto 0);  -- pio_captura_2_s1_translator:uav_readdata -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                  : std_logic;                      -- pio_captura_2_s1_translator:uav_readdatavalid -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                    : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_captura_2_s1_translator:uav_debugaccess
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                     : std_logic_vector(3 downto 0);   -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_captura_2_s1_translator:uav_byteenable
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket             : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                   : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket           : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data                    : std_logic_vector(104 downto 0); -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                   : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket          : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket        : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                 : std_logic_vector(104 downto 0); -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid              : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data               : std_logic_vector(33 downto 0);  -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready              : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                    : std_logic;                      -- pio_captura_3_s1_translator:uav_waitrequest -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                     : std_logic_vector(2 downto 0);   -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_captura_3_s1_translator:uav_burstcount
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata                      : std_logic_vector(31 downto 0);  -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_captura_3_s1_translator:uav_writedata
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_address                        : std_logic_vector(24 downto 0);  -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_captura_3_s1_translator:uav_address
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_write                          : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_captura_3_s1_translator:uav_write
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_lock                           : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_captura_3_s1_translator:uav_lock
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_read                           : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_captura_3_s1_translator:uav_read
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata                       : std_logic_vector(31 downto 0);  -- pio_captura_3_s1_translator:uav_readdata -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                  : std_logic;                      -- pio_captura_3_s1_translator:uav_readdatavalid -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                    : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_captura_3_s1_translator:uav_debugaccess
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                     : std_logic_vector(3 downto 0);   -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_captura_3_s1_translator:uav_byteenable
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket             : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                   : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket           : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data                    : std_logic_vector(104 downto 0); -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                   : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket          : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket        : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                 : std_logic_vector(104 downto 0); -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid              : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data               : std_logic_vector(33 downto 0);  -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready              : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                    : std_logic;                      -- pio_captura_4_s1_translator:uav_waitrequest -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                     : std_logic_vector(2 downto 0);   -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_captura_4_s1_translator:uav_burstcount
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata                      : std_logic_vector(31 downto 0);  -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_captura_4_s1_translator:uav_writedata
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_address                        : std_logic_vector(24 downto 0);  -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_captura_4_s1_translator:uav_address
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_write                          : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_captura_4_s1_translator:uav_write
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_lock                           : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_captura_4_s1_translator:uav_lock
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_read                           : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_captura_4_s1_translator:uav_read
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata                       : std_logic_vector(31 downto 0);  -- pio_captura_4_s1_translator:uav_readdata -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                  : std_logic;                      -- pio_captura_4_s1_translator:uav_readdatavalid -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                    : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_captura_4_s1_translator:uav_debugaccess
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                     : std_logic_vector(3 downto 0);   -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_captura_4_s1_translator:uav_byteenable
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket             : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                   : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket           : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data                    : std_logic_vector(104 downto 0); -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                   : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket          : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket        : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                 : std_logic_vector(104 downto 0); -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid              : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data               : std_logic_vector(33 downto 0);  -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready              : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                        : std_logic;                      -- pio_in_32_s1_translator:uav_waitrequest -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                         : std_logic_vector(2 downto 0);   -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_in_32_s1_translator:uav_burstcount
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_writedata                          : std_logic_vector(31 downto 0);  -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_in_32_s1_translator:uav_writedata
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_address                            : std_logic_vector(24 downto 0);  -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_in_32_s1_translator:uav_address
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_write                              : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_in_32_s1_translator:uav_write
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_lock                               : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_in_32_s1_translator:uav_lock
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_read                               : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_in_32_s1_translator:uav_read
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_readdata                           : std_logic_vector(31 downto 0);  -- pio_in_32_s1_translator:uav_readdata -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                      : std_logic;                      -- pio_in_32_s1_translator:uav_readdatavalid -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                        : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_in_32_s1_translator:uav_debugaccess
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                         : std_logic_vector(3 downto 0);   -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_in_32_s1_translator:uav_byteenable
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                 : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                       : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket               : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rf_source_data                        : std_logic_vector(104 downto 0); -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                       : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket              : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                    : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket            : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                     : std_logic_vector(104 downto 0); -- pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                    : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                  : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                   : std_logic_vector(33 downto 0);  -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                  : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                   : std_logic;                      -- lcd_control_slave_translator:uav_waitrequest -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                    : std_logic_vector(2 downto 0);   -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_control_slave_translator:uav_burstcount
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                     : std_logic_vector(31 downto 0);  -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_control_slave_translator:uav_writedata
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address                       : std_logic_vector(24 downto 0);  -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> lcd_control_slave_translator:uav_address
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write                         : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> lcd_control_slave_translator:uav_write
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                          : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_control_slave_translator:uav_lock
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read                          : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> lcd_control_slave_translator:uav_read
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                      : std_logic_vector(31 downto 0);  -- lcd_control_slave_translator:uav_readdata -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                 : std_logic;                      -- lcd_control_slave_translator:uav_readdatavalid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                   : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_control_slave_translator:uav_debugaccess
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                    : std_logic_vector(3 downto 0);   -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_control_slave_translator:uav_byteenable
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket            : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                  : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket          : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                   : std_logic_vector(104 downto 0); -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                  : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket         : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid               : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket       : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                : std_logic_vector(104 downto 0); -- lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready               : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid             : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data              : std_logic_vector(33 downto 0);  -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready             : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest              : std_logic;                      -- DM9000A_avalon_slave_0_translator:uav_waitrequest -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount               : std_logic_vector(2 downto 0);   -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> DM9000A_avalon_slave_0_translator:uav_burstcount
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata                : std_logic_vector(31 downto 0);  -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> DM9000A_avalon_slave_0_translator:uav_writedata
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                  : std_logic_vector(24 downto 0);  -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> DM9000A_avalon_slave_0_translator:uav_address
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                    : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> DM9000A_avalon_slave_0_translator:uav_write
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                     : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> DM9000A_avalon_slave_0_translator:uav_lock
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                     : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> DM9000A_avalon_slave_0_translator:uav_read
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                 : std_logic_vector(31 downto 0);  -- DM9000A_avalon_slave_0_translator:uav_readdata -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid            : std_logic;                      -- DM9000A_avalon_slave_0_translator:uav_readdatavalid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess              : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> DM9000A_avalon_slave_0_translator:uav_debugaccess
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable               : std_logic_vector(3 downto 0);   -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> DM9000A_avalon_slave_0_translator:uav_byteenable
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket       : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid             : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket     : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data              : std_logic_vector(104 downto 0); -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready             : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid          : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket  : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data           : std_logic_vector(104 downto 0); -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready          : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid        : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         : std_logic_vector(33 downto 0);  -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready        : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket             : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                   : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket           : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data                    : std_logic_vector(103 downto 0); -- cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                   : std_logic;                      -- addr_router:sink_ready -> cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                    : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid                          : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                  : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_data                           : std_logic_vector(103 downto 0); -- cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready                          : std_logic;                      -- addr_router_001:sink_ready -> cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket               : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                     : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket             : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                      : std_logic_vector(103 downto 0); -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                     : std_logic;                      -- id_router:sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                            : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid                                  : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                          : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_data                                   : std_logic_vector(85 downto 0);  -- sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready                                  : std_logic;                      -- id_router_001:sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(103 downto 0); -- system_id_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal system_id_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                      -- id_router_002:sink_ready -> system_id_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                       : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid                             : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                     : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data                              : std_logic_vector(103 downto 0); -- pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready                             : std_logic;                      -- id_router_003:sink_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket              : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                    : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket            : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                     : std_logic_vector(103 downto 0); -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                    : std_logic;                      -- id_router_004:sink_ready -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                          : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                                : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                        : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data                                 : std_logic_vector(103 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                                : std_logic;                      -- id_router_005:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                          : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid                                : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                        : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data                                 : std_logic_vector(103 downto 0); -- timer_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready                                : std_logic;                      -- id_router_006:sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                        : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rp_valid                              : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                      : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rp_data                               : std_logic_vector(103 downto 0); -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rp_ready                              : std_logic;                      -- id_router_007:sink_ready -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                  : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rp_valid                        : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rp_data                         : std_logic_vector(103 downto 0); -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	signal pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rp_ready                        : std_logic;                      -- id_router_008:sink_ready -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                       : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rp_valid                             : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                     : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rp_data                              : std_logic_vector(103 downto 0); -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	signal pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rp_ready                             : std_logic;                      -- id_router_009:sink_ready -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                      : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rp_valid                            : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                    : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rp_data                             : std_logic_vector(103 downto 0); -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	signal pio_out_red_s1_translator_avalon_universal_slave_0_agent_rp_ready                            : std_logic;                      -- id_router_010:sink_ready -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                    : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rp_valid                          : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                  : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rp_data                           : std_logic_vector(103 downto 0); -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	signal pio_out_green_s1_translator_avalon_universal_slave_0_agent_rp_ready                          : std_logic;                      -- id_router_011:sink_ready -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                      : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rp_valid                            : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                    : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rp_data                             : std_logic_vector(103 downto 0); -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	signal pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rp_ready                            : std_logic;                      -- id_router_012:sink_ready -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                  : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rp_valid                        : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rp_data                         : std_logic_vector(103 downto 0); -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	signal pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rp_ready                        : std_logic;                      -- id_router_013:sink_ready -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                       : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rp_valid                             : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                     : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rp_data                              : std_logic_vector(103 downto 0); -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	signal pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rp_ready                             : std_logic;                      -- id_router_014:sink_ready -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                        : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rp_valid                              : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                      : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rp_data                               : std_logic_vector(103 downto 0); -- pio_direc_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	signal pio_direc_s1_translator_avalon_universal_slave_0_agent_rp_ready                              : std_logic;                      -- id_router_015:sink_ready -> pio_direc_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                    : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid                          : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                  : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rp_data                           : std_logic_vector(103 downto 0); -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	signal pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready                          : std_logic;                      -- id_router_016:sink_ready -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                           : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rp_valid                                 : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                         : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rp_data                                  : std_logic_vector(103 downto 0); -- pio_wr_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	signal pio_wr_s1_translator_avalon_universal_slave_0_agent_rp_ready                                 : std_logic;                      -- id_router_017:sink_ready -> pio_wr_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                   : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rp_valid                         : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                 : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rp_data                          : std_logic_vector(103 downto 0); -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	signal pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rp_ready                         : std_logic;                      -- id_router_018:sink_ready -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                        : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rp_valid                              : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                      : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rp_data                               : std_logic_vector(103 downto 0); -- pio_datos_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	signal pio_datos_s1_translator_avalon_universal_slave_0_agent_rp_ready                              : std_logic;                      -- id_router_019:sink_ready -> pio_datos_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                      : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket              : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rp_data                       : std_logic_vector(103 downto 0); -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	signal pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                      : std_logic;                      -- id_router_020:sink_ready -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rp_valid                      : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket              : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rp_data                       : std_logic_vector(103 downto 0); -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	signal pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rp_ready                      : std_logic;                      -- id_router_021:sink_ready -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rp_valid                      : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket              : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rp_data                       : std_logic_vector(103 downto 0); -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	signal pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rp_ready                      : std_logic;                      -- id_router_022:sink_ready -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_023:sink_endofpacket
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rp_valid                      : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_023:sink_valid
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket              : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_023:sink_startofpacket
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rp_data                       : std_logic_vector(103 downto 0); -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_023:sink_data
	signal pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rp_ready                      : std_logic;                      -- id_router_023:sink_ready -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_024:sink_endofpacket
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rp_valid                      : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_024:sink_valid
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket              : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_024:sink_startofpacket
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rp_data                       : std_logic_vector(103 downto 0); -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_024:sink_data
	signal pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rp_ready                      : std_logic;                      -- id_router_024:sink_ready -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                    : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_025:sink_endofpacket
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                          : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_025:sink_valid
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                  : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_025:sink_startofpacket
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rp_data                           : std_logic_vector(103 downto 0); -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_025:sink_data
	signal pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                          : std_logic;                      -- id_router_025:sink_ready -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                    : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_026:sink_endofpacket
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rp_valid                          : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_026:sink_valid
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                  : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_026:sink_startofpacket
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rp_data                           : std_logic_vector(103 downto 0); -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_026:sink_data
	signal pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rp_ready                          : std_logic;                      -- id_router_026:sink_ready -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                    : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_027:sink_endofpacket
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rp_valid                          : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_027:sink_valid
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                  : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_027:sink_startofpacket
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rp_data                           : std_logic_vector(103 downto 0); -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_027:sink_data
	signal pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rp_ready                          : std_logic;                      -- id_router_027:sink_ready -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                    : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_028:sink_endofpacket
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rp_valid                          : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_028:sink_valid
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                  : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_028:sink_startofpacket
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rp_data                           : std_logic_vector(103 downto 0); -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_028:sink_data
	signal pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rp_ready                          : std_logic;                      -- id_router_028:sink_ready -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                    : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_029:sink_endofpacket
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rp_valid                          : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_029:sink_valid
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                  : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_029:sink_startofpacket
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rp_data                           : std_logic_vector(103 downto 0); -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_029:sink_data
	signal pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rp_ready                          : std_logic;                      -- id_router_029:sink_ready -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                        : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_030:sink_endofpacket
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rp_valid                              : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_030:sink_valid
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                      : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_030:sink_startofpacket
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rp_data                               : std_logic_vector(103 downto 0); -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_030:sink_data
	signal pio_in_32_s1_translator_avalon_universal_slave_0_agent_rp_ready                              : std_logic;                      -- id_router_030:sink_ready -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                   : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_031:sink_endofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                         : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_031:sink_valid
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                 : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_031:sink_startofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data                          : std_logic_vector(103 downto 0); -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_031:sink_data
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                         : std_logic;                      -- id_router_031:sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket              : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_032:sink_endofpacket
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                    : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_032:sink_valid
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket            : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_032:sink_startofpacket
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                     : std_logic_vector(103 downto 0); -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_032:sink_data
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                    : std_logic;                      -- id_router_032:sink_ready -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal addr_router_src_endofpacket                                                                  : std_logic;                      -- addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	signal addr_router_src_valid                                                                        : std_logic;                      -- addr_router:src_valid -> limiter:cmd_sink_valid
	signal addr_router_src_startofpacket                                                                : std_logic;                      -- addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	signal addr_router_src_data                                                                         : std_logic_vector(103 downto 0); -- addr_router:src_data -> limiter:cmd_sink_data
	signal addr_router_src_channel                                                                      : std_logic_vector(32 downto 0);  -- addr_router:src_channel -> limiter:cmd_sink_channel
	signal addr_router_src_ready                                                                        : std_logic;                      -- limiter:cmd_sink_ready -> addr_router:src_ready
	signal limiter_rsp_src_endofpacket                                                                  : std_logic;                      -- limiter:rsp_src_endofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_rsp_src_valid                                                                        : std_logic;                      -- limiter:rsp_src_valid -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_rsp_src_startofpacket                                                                : std_logic;                      -- limiter:rsp_src_startofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_rsp_src_data                                                                         : std_logic_vector(103 downto 0); -- limiter:rsp_src_data -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_rsp_src_channel                                                                      : std_logic_vector(32 downto 0);  -- limiter:rsp_src_channel -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_rsp_src_ready                                                                        : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	signal burst_adapter_source0_endofpacket                                                            : std_logic;                      -- burst_adapter:source0_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_source0_valid                                                                  : std_logic;                      -- burst_adapter:source0_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_source0_startofpacket                                                          : std_logic;                      -- burst_adapter:source0_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_source0_data                                                                   : std_logic_vector(85 downto 0);  -- burst_adapter:source0_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_source0_ready                                                                  : std_logic;                      -- sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	signal burst_adapter_source0_channel                                                                : std_logic_vector(32 downto 0);  -- burst_adapter:source0_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal rst_controller_reset_out_reset                                                               : std_logic;                      -- rst_controller:reset_out -> [DM9000A_avalon_slave_0_translator:reset, DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, burst_adapter:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cpu_data_master_translator:reset, cpu_data_master_translator_avalon_universal_master_0_agent:reset, cpu_instruction_master_translator:reset, cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_jtag_debug_module_translator:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:in_reset, crosser_001:out_reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, id_router_020:reset, id_router_021:reset, id_router_022:reset, id_router_023:reset, id_router_024:reset, id_router_025:reset, id_router_026:reset, id_router_027:reset, id_router_028:reset, id_router_029:reset, id_router_030:reset, id_router_031:reset, id_router_032:reset, irq_mapper:reset, lcd_control_slave_translator:reset, lcd_control_slave_translator_avalon_universal_slave_0_agent:reset, lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, pio_async_reset_s1_translator:reset, pio_async_reset_s1_translator_avalon_universal_slave_0_agent:reset, pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_captura_0_s1_translator:reset, pio_captura_0_s1_translator_avalon_universal_slave_0_agent:reset, pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_captura_1_s1_translator:reset, pio_captura_1_s1_translator_avalon_universal_slave_0_agent:reset, pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_captura_2_s1_translator:reset, pio_captura_2_s1_translator_avalon_universal_slave_0_agent:reset, pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_captura_3_s1_translator:reset, pio_captura_3_s1_translator_avalon_universal_slave_0_agent:reset, pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_captura_4_s1_translator:reset, pio_captura_4_s1_translator_avalon_universal_slave_0_agent:reset, pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_compara_int_0_s1_translator:reset, pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:reset, pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_compara_int_1_s1_translator:reset, pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:reset, pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_compara_int_2_s1_translator:reset, pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:reset, pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_compara_int_3_s1_translator:reset, pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:reset, pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_compara_int_4_s1_translator:reset, pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:reset, pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_datos_s1_translator:reset, pio_datos_s1_translator_avalon_universal_slave_0_agent:reset, pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_direc_ram_s1_translator:reset, pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:reset, pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_direc_s1_translator:reset, pio_direc_s1_translator_avalon_universal_slave_0_agent:reset, pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_en_mux_s1_translator:reset, pio_en_mux_s1_translator_avalon_universal_slave_0_agent:reset, pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_in_32_s1_translator:reset, pio_in_32_s1_translator_avalon_universal_slave_0_agent:reset, pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_in_ext_s1_translator:reset, pio_in_ext_s1_translator_avalon_universal_slave_0_agent:reset, pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_in_key_edge_s1_translator:reset, pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:reset, pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_in_sw_s1_translator:reset, pio_in_sw_s1_translator_avalon_universal_slave_0_agent:reset, pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_out_ext_s1_translator:reset, pio_out_ext_s1_translator_avalon_universal_slave_0_agent:reset, pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_out_green_s1_translator:reset, pio_out_green_s1_translator_avalon_universal_slave_0_agent:reset, pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_out_red_s1_translator:reset, pio_out_red_s1_translator_avalon_universal_slave_0_agent:reset, pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_sel_salida_s1_translator:reset, pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:reset, pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_wr_s1_translator:reset, pio_wr_s1_translator_avalon_universal_slave_0_agent:reset, pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_022:reset, rsp_xbar_demux_023:reset, rsp_xbar_demux_024:reset, rsp_xbar_demux_025:reset, rsp_xbar_demux_026:reset, rsp_xbar_demux_027:reset, rsp_xbar_demux_028:reset, rsp_xbar_demux_029:reset, rsp_xbar_demux_030:reset, rsp_xbar_demux_031:reset, rsp_xbar_demux_032:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_reset_out_reset:in, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, system_id_control_slave_translator:reset, system_id_control_slave_translator_avalon_universal_slave_0_agent:reset, system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_1_s1_translator:reset, timer_1_s1_translator_avalon_universal_slave_0_agent:reset, timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, uart_avalon_jtag_slave_translator:reset, uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset]
	signal rst_controller_001_reset_out_reset                                                           : std_logic;                      -- rst_controller_001:reset_out -> [crosser:out_reset, crosser_001:in_reset, id_router_003:reset, pll:reset, pll_pll_slave_translator:reset, pll_pll_slave_translator_avalon_universal_slave_0_agent:reset, pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_003:reset]
	signal cmd_xbar_demux_src0_endofpacket                                                              : std_logic;                      -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                    : std_logic;                      -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                            : std_logic;                      -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                     : std_logic_vector(103 downto 0); -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                  : std_logic_vector(32 downto 0);  -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                    : std_logic;                      -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                              : std_logic;                      -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                    : std_logic;                      -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                            : std_logic;                      -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                     : std_logic_vector(103 downto 0); -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                  : std_logic_vector(32 downto 0);  -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                    : std_logic;                      -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_src2_endofpacket                                                              : std_logic;                      -- cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	signal cmd_xbar_demux_src2_valid                                                                    : std_logic;                      -- cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	signal cmd_xbar_demux_src2_startofpacket                                                            : std_logic;                      -- cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	signal cmd_xbar_demux_src2_data                                                                     : std_logic_vector(103 downto 0); -- cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	signal cmd_xbar_demux_src2_channel                                                                  : std_logic_vector(32 downto 0);  -- cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	signal cmd_xbar_demux_src2_ready                                                                    : std_logic;                      -- cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                          : std_logic;                      -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                : std_logic;                      -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                        : std_logic;                      -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                 : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                              : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                : std_logic;                      -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                          : std_logic;                      -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                : std_logic;                      -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                        : std_logic;                      -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                 : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                              : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                : std_logic;                      -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src2_endofpacket                                                          : std_logic;                      -- cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                                : std_logic;                      -- cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                        : std_logic;                      -- cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                                 : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	signal cmd_xbar_demux_001_src2_channel                                                              : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	signal cmd_xbar_demux_001_src2_ready                                                                : std_logic;                      -- cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	signal cmd_xbar_demux_001_src4_endofpacket                                                          : std_logic;                      -- cmd_xbar_demux_001:src4_endofpacket -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src4_valid                                                                : std_logic;                      -- cmd_xbar_demux_001:src4_valid -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src4_startofpacket                                                        : std_logic;                      -- cmd_xbar_demux_001:src4_startofpacket -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src4_data                                                                 : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src4_data -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src4_channel                                                              : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src4_channel -> uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src5_endofpacket                                                          : std_logic;                      -- cmd_xbar_demux_001:src5_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src5_valid                                                                : std_logic;                      -- cmd_xbar_demux_001:src5_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src5_startofpacket                                                        : std_logic;                      -- cmd_xbar_demux_001:src5_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src5_data                                                                 : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src5_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src5_channel                                                              : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src5_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src6_endofpacket                                                          : std_logic;                      -- cmd_xbar_demux_001:src6_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src6_valid                                                                : std_logic;                      -- cmd_xbar_demux_001:src6_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src6_startofpacket                                                        : std_logic;                      -- cmd_xbar_demux_001:src6_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src6_data                                                                 : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src6_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src6_channel                                                              : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src6_channel -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src7_endofpacket                                                          : std_logic;                      -- cmd_xbar_demux_001:src7_endofpacket -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src7_valid                                                                : std_logic;                      -- cmd_xbar_demux_001:src7_valid -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src7_startofpacket                                                        : std_logic;                      -- cmd_xbar_demux_001:src7_startofpacket -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src7_data                                                                 : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src7_data -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src7_channel                                                              : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src7_channel -> pio_in_sw_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src8_endofpacket                                                          : std_logic;                      -- cmd_xbar_demux_001:src8_endofpacket -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src8_valid                                                                : std_logic;                      -- cmd_xbar_demux_001:src8_valid -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src8_startofpacket                                                        : std_logic;                      -- cmd_xbar_demux_001:src8_startofpacket -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src8_data                                                                 : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src8_data -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src8_channel                                                              : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src8_channel -> pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src9_endofpacket                                                          : std_logic;                      -- cmd_xbar_demux_001:src9_endofpacket -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src9_valid                                                                : std_logic;                      -- cmd_xbar_demux_001:src9_valid -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src9_startofpacket                                                        : std_logic;                      -- cmd_xbar_demux_001:src9_startofpacket -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src9_data                                                                 : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src9_data -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src9_channel                                                              : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src9_channel -> pio_in_ext_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src10_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src10_endofpacket -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src10_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src10_valid -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src10_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src10_startofpacket -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src10_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src10_data -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src10_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src10_channel -> pio_out_red_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src11_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src11_endofpacket -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src11_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src11_valid -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src11_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src11_startofpacket -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src11_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src11_data -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src11_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src11_channel -> pio_out_green_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src12_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src12_endofpacket -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src12_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src12_valid -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src12_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src12_startofpacket -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src12_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src12_data -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src12_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src12_channel -> pio_out_ext_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src13_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src13_endofpacket -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src13_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src13_valid -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src13_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src13_startofpacket -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src13_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src13_data -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src13_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src13_channel -> pio_async_reset_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src14_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src14_endofpacket -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src14_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src14_valid -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src14_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src14_startofpacket -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src14_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src14_data -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src14_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src14_channel -> pio_en_mux_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src15_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src15_endofpacket -> pio_direc_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src15_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src15_valid -> pio_direc_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src15_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src15_startofpacket -> pio_direc_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src15_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src15_data -> pio_direc_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src15_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src15_channel -> pio_direc_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src16_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src16_endofpacket -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src16_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src16_valid -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src16_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src16_startofpacket -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src16_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src16_data -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src16_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src16_channel -> pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src17_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src17_endofpacket -> pio_wr_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src17_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src17_valid -> pio_wr_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src17_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src17_startofpacket -> pio_wr_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src17_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src17_data -> pio_wr_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src17_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src17_channel -> pio_wr_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src18_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src18_endofpacket -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src18_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src18_valid -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src18_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src18_startofpacket -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src18_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src18_data -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src18_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src18_channel -> pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src19_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src19_endofpacket -> pio_datos_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src19_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src19_valid -> pio_datos_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src19_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src19_startofpacket -> pio_datos_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src19_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src19_data -> pio_datos_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src19_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src19_channel -> pio_datos_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src20_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src20_endofpacket -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src20_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src20_valid -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src20_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src20_startofpacket -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src20_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src20_data -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src20_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src20_channel -> pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src21_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src21_endofpacket -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src21_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src21_valid -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src21_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src21_startofpacket -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src21_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src21_data -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src21_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src21_channel -> pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src22_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src22_endofpacket -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src22_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src22_valid -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src22_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src22_startofpacket -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src22_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src22_data -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src22_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src22_channel -> pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src23_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src23_endofpacket -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src23_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src23_valid -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src23_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src23_startofpacket -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src23_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src23_data -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src23_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src23_channel -> pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src24_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src24_endofpacket -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src24_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src24_valid -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src24_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src24_startofpacket -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src24_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src24_data -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src24_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src24_channel -> pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src25_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src25_endofpacket -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src25_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src25_valid -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src25_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src25_startofpacket -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src25_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src25_data -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src25_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src25_channel -> pio_captura_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src26_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src26_endofpacket -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src26_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src26_valid -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src26_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src26_startofpacket -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src26_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src26_data -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src26_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src26_channel -> pio_captura_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src27_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src27_endofpacket -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src27_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src27_valid -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src27_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src27_startofpacket -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src27_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src27_data -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src27_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src27_channel -> pio_captura_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src28_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src28_endofpacket -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src28_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src28_valid -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src28_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src28_startofpacket -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src28_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src28_data -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src28_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src28_channel -> pio_captura_3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src29_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src29_endofpacket -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src29_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src29_valid -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src29_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src29_startofpacket -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src29_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src29_data -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src29_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src29_channel -> pio_captura_4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src30_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src30_endofpacket -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src30_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src30_valid -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src30_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src30_startofpacket -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src30_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src30_data -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src30_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src30_channel -> pio_in_32_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src31_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src31_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src31_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src31_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src31_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src31_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src31_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src31_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src31_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src31_channel -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src32_endofpacket                                                         : std_logic;                      -- cmd_xbar_demux_001:src32_endofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src32_valid                                                               : std_logic;                      -- cmd_xbar_demux_001:src32_valid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src32_startofpacket                                                       : std_logic;                      -- cmd_xbar_demux_001:src32_startofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src32_data                                                                : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src32_data -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src32_channel                                                             : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src32_channel -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal rsp_xbar_demux_src0_endofpacket                                                              : std_logic;                      -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                    : std_logic;                      -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                            : std_logic;                      -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                     : std_logic_vector(103 downto 0); -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                  : std_logic_vector(32 downto 0);  -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                    : std_logic;                      -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                              : std_logic;                      -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                    : std_logic;                      -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                            : std_logic;                      -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                     : std_logic_vector(103 downto 0); -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                  : std_logic_vector(32 downto 0);  -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                    : std_logic;                      -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                : std_logic;                      -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_002_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_002_src1_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal rsp_xbar_demux_002_src1_valid                                                                : std_logic;                      -- rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	signal rsp_xbar_demux_002_src1_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal rsp_xbar_demux_002_src1_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	signal rsp_xbar_demux_002_src1_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_002_src1_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	signal rsp_xbar_demux_004_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	signal rsp_xbar_demux_004_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	signal rsp_xbar_demux_005_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	signal rsp_xbar_demux_005_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	signal rsp_xbar_demux_005_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	signal rsp_xbar_demux_006_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	signal rsp_xbar_demux_006_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	signal rsp_xbar_demux_007_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	signal rsp_xbar_demux_007_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	signal rsp_xbar_demux_008_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	signal rsp_xbar_demux_008_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	signal rsp_xbar_demux_008_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	signal rsp_xbar_demux_008_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	signal rsp_xbar_demux_008_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	signal rsp_xbar_demux_008_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	signal rsp_xbar_demux_009_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	signal rsp_xbar_demux_009_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	signal rsp_xbar_demux_009_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	signal rsp_xbar_demux_009_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	signal rsp_xbar_demux_009_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	signal rsp_xbar_demux_009_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	signal rsp_xbar_demux_010_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	signal rsp_xbar_demux_010_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	signal rsp_xbar_demux_010_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	signal rsp_xbar_demux_010_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	signal rsp_xbar_demux_010_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	signal rsp_xbar_demux_010_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	signal rsp_xbar_demux_011_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	signal rsp_xbar_demux_011_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	signal rsp_xbar_demux_011_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	signal rsp_xbar_demux_011_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	signal rsp_xbar_demux_011_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	signal rsp_xbar_demux_011_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	signal rsp_xbar_demux_012_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	signal rsp_xbar_demux_012_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	signal rsp_xbar_demux_012_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	signal rsp_xbar_demux_012_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	signal rsp_xbar_demux_012_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	signal rsp_xbar_demux_012_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	signal rsp_xbar_demux_013_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	signal rsp_xbar_demux_013_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	signal rsp_xbar_demux_013_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	signal rsp_xbar_demux_013_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	signal rsp_xbar_demux_013_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	signal rsp_xbar_demux_013_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	signal rsp_xbar_demux_014_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	signal rsp_xbar_demux_014_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink14_valid
	signal rsp_xbar_demux_014_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	signal rsp_xbar_demux_014_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink14_data
	signal rsp_xbar_demux_014_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink14_channel
	signal rsp_xbar_demux_014_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src0_ready
	signal rsp_xbar_demux_015_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	signal rsp_xbar_demux_015_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	signal rsp_xbar_demux_015_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	signal rsp_xbar_demux_015_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	signal rsp_xbar_demux_015_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	signal rsp_xbar_demux_015_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	signal rsp_xbar_demux_016_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	signal rsp_xbar_demux_016_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_001:sink16_valid
	signal rsp_xbar_demux_016_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	signal rsp_xbar_demux_016_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_001:sink16_data
	signal rsp_xbar_demux_016_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_001:sink16_channel
	signal rsp_xbar_demux_016_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src0_ready
	signal rsp_xbar_demux_017_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	signal rsp_xbar_demux_017_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_001:sink17_valid
	signal rsp_xbar_demux_017_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	signal rsp_xbar_demux_017_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_001:sink17_data
	signal rsp_xbar_demux_017_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_001:sink17_channel
	signal rsp_xbar_demux_017_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink17_ready -> rsp_xbar_demux_017:src0_ready
	signal rsp_xbar_demux_018_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	signal rsp_xbar_demux_018_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_001:sink18_valid
	signal rsp_xbar_demux_018_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	signal rsp_xbar_demux_018_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_001:sink18_data
	signal rsp_xbar_demux_018_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_001:sink18_channel
	signal rsp_xbar_demux_018_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink18_ready -> rsp_xbar_demux_018:src0_ready
	signal rsp_xbar_demux_019_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_001:sink19_endofpacket
	signal rsp_xbar_demux_019_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_001:sink19_valid
	signal rsp_xbar_demux_019_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_001:sink19_startofpacket
	signal rsp_xbar_demux_019_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_001:sink19_data
	signal rsp_xbar_demux_019_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_001:sink19_channel
	signal rsp_xbar_demux_019_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink19_ready -> rsp_xbar_demux_019:src0_ready
	signal rsp_xbar_demux_020_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux_001:sink20_endofpacket
	signal rsp_xbar_demux_020_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux_001:sink20_valid
	signal rsp_xbar_demux_020_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux_001:sink20_startofpacket
	signal rsp_xbar_demux_020_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_020:src0_data -> rsp_xbar_mux_001:sink20_data
	signal rsp_xbar_demux_020_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux_001:sink20_channel
	signal rsp_xbar_demux_020_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink20_ready -> rsp_xbar_demux_020:src0_ready
	signal rsp_xbar_demux_021_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux_001:sink21_endofpacket
	signal rsp_xbar_demux_021_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux_001:sink21_valid
	signal rsp_xbar_demux_021_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux_001:sink21_startofpacket
	signal rsp_xbar_demux_021_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_021:src0_data -> rsp_xbar_mux_001:sink21_data
	signal rsp_xbar_demux_021_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux_001:sink21_channel
	signal rsp_xbar_demux_021_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink21_ready -> rsp_xbar_demux_021:src0_ready
	signal rsp_xbar_demux_022_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux_001:sink22_endofpacket
	signal rsp_xbar_demux_022_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux_001:sink22_valid
	signal rsp_xbar_demux_022_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux_001:sink22_startofpacket
	signal rsp_xbar_demux_022_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_022:src0_data -> rsp_xbar_mux_001:sink22_data
	signal rsp_xbar_demux_022_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux_001:sink22_channel
	signal rsp_xbar_demux_022_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink22_ready -> rsp_xbar_demux_022:src0_ready
	signal rsp_xbar_demux_023_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_023:src0_endofpacket -> rsp_xbar_mux_001:sink23_endofpacket
	signal rsp_xbar_demux_023_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_023:src0_valid -> rsp_xbar_mux_001:sink23_valid
	signal rsp_xbar_demux_023_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_023:src0_startofpacket -> rsp_xbar_mux_001:sink23_startofpacket
	signal rsp_xbar_demux_023_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_023:src0_data -> rsp_xbar_mux_001:sink23_data
	signal rsp_xbar_demux_023_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_023:src0_channel -> rsp_xbar_mux_001:sink23_channel
	signal rsp_xbar_demux_023_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink23_ready -> rsp_xbar_demux_023:src0_ready
	signal rsp_xbar_demux_024_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_024:src0_endofpacket -> rsp_xbar_mux_001:sink24_endofpacket
	signal rsp_xbar_demux_024_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_024:src0_valid -> rsp_xbar_mux_001:sink24_valid
	signal rsp_xbar_demux_024_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_024:src0_startofpacket -> rsp_xbar_mux_001:sink24_startofpacket
	signal rsp_xbar_demux_024_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_024:src0_data -> rsp_xbar_mux_001:sink24_data
	signal rsp_xbar_demux_024_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_024:src0_channel -> rsp_xbar_mux_001:sink24_channel
	signal rsp_xbar_demux_024_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink24_ready -> rsp_xbar_demux_024:src0_ready
	signal rsp_xbar_demux_025_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_025:src0_endofpacket -> rsp_xbar_mux_001:sink25_endofpacket
	signal rsp_xbar_demux_025_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_025:src0_valid -> rsp_xbar_mux_001:sink25_valid
	signal rsp_xbar_demux_025_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_025:src0_startofpacket -> rsp_xbar_mux_001:sink25_startofpacket
	signal rsp_xbar_demux_025_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_025:src0_data -> rsp_xbar_mux_001:sink25_data
	signal rsp_xbar_demux_025_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_025:src0_channel -> rsp_xbar_mux_001:sink25_channel
	signal rsp_xbar_demux_025_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink25_ready -> rsp_xbar_demux_025:src0_ready
	signal rsp_xbar_demux_026_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_026:src0_endofpacket -> rsp_xbar_mux_001:sink26_endofpacket
	signal rsp_xbar_demux_026_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_026:src0_valid -> rsp_xbar_mux_001:sink26_valid
	signal rsp_xbar_demux_026_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_026:src0_startofpacket -> rsp_xbar_mux_001:sink26_startofpacket
	signal rsp_xbar_demux_026_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_026:src0_data -> rsp_xbar_mux_001:sink26_data
	signal rsp_xbar_demux_026_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_026:src0_channel -> rsp_xbar_mux_001:sink26_channel
	signal rsp_xbar_demux_026_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink26_ready -> rsp_xbar_demux_026:src0_ready
	signal rsp_xbar_demux_027_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_027:src0_endofpacket -> rsp_xbar_mux_001:sink27_endofpacket
	signal rsp_xbar_demux_027_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_027:src0_valid -> rsp_xbar_mux_001:sink27_valid
	signal rsp_xbar_demux_027_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_027:src0_startofpacket -> rsp_xbar_mux_001:sink27_startofpacket
	signal rsp_xbar_demux_027_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_027:src0_data -> rsp_xbar_mux_001:sink27_data
	signal rsp_xbar_demux_027_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_027:src0_channel -> rsp_xbar_mux_001:sink27_channel
	signal rsp_xbar_demux_027_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink27_ready -> rsp_xbar_demux_027:src0_ready
	signal rsp_xbar_demux_028_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_028:src0_endofpacket -> rsp_xbar_mux_001:sink28_endofpacket
	signal rsp_xbar_demux_028_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_028:src0_valid -> rsp_xbar_mux_001:sink28_valid
	signal rsp_xbar_demux_028_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_028:src0_startofpacket -> rsp_xbar_mux_001:sink28_startofpacket
	signal rsp_xbar_demux_028_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_028:src0_data -> rsp_xbar_mux_001:sink28_data
	signal rsp_xbar_demux_028_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_028:src0_channel -> rsp_xbar_mux_001:sink28_channel
	signal rsp_xbar_demux_028_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink28_ready -> rsp_xbar_demux_028:src0_ready
	signal rsp_xbar_demux_029_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_029:src0_endofpacket -> rsp_xbar_mux_001:sink29_endofpacket
	signal rsp_xbar_demux_029_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_029:src0_valid -> rsp_xbar_mux_001:sink29_valid
	signal rsp_xbar_demux_029_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_029:src0_startofpacket -> rsp_xbar_mux_001:sink29_startofpacket
	signal rsp_xbar_demux_029_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_029:src0_data -> rsp_xbar_mux_001:sink29_data
	signal rsp_xbar_demux_029_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_029:src0_channel -> rsp_xbar_mux_001:sink29_channel
	signal rsp_xbar_demux_029_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink29_ready -> rsp_xbar_demux_029:src0_ready
	signal rsp_xbar_demux_030_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_030:src0_endofpacket -> rsp_xbar_mux_001:sink30_endofpacket
	signal rsp_xbar_demux_030_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_030:src0_valid -> rsp_xbar_mux_001:sink30_valid
	signal rsp_xbar_demux_030_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_030:src0_startofpacket -> rsp_xbar_mux_001:sink30_startofpacket
	signal rsp_xbar_demux_030_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_030:src0_data -> rsp_xbar_mux_001:sink30_data
	signal rsp_xbar_demux_030_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_030:src0_channel -> rsp_xbar_mux_001:sink30_channel
	signal rsp_xbar_demux_030_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink30_ready -> rsp_xbar_demux_030:src0_ready
	signal rsp_xbar_demux_031_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_031:src0_endofpacket -> rsp_xbar_mux_001:sink31_endofpacket
	signal rsp_xbar_demux_031_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_031:src0_valid -> rsp_xbar_mux_001:sink31_valid
	signal rsp_xbar_demux_031_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_031:src0_startofpacket -> rsp_xbar_mux_001:sink31_startofpacket
	signal rsp_xbar_demux_031_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_031:src0_data -> rsp_xbar_mux_001:sink31_data
	signal rsp_xbar_demux_031_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_031:src0_channel -> rsp_xbar_mux_001:sink31_channel
	signal rsp_xbar_demux_031_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink31_ready -> rsp_xbar_demux_031:src0_ready
	signal rsp_xbar_demux_032_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_032:src0_endofpacket -> rsp_xbar_mux_001:sink32_endofpacket
	signal rsp_xbar_demux_032_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_032:src0_valid -> rsp_xbar_mux_001:sink32_valid
	signal rsp_xbar_demux_032_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_032:src0_startofpacket -> rsp_xbar_mux_001:sink32_startofpacket
	signal rsp_xbar_demux_032_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_032:src0_data -> rsp_xbar_mux_001:sink32_data
	signal rsp_xbar_demux_032_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_032:src0_channel -> rsp_xbar_mux_001:sink32_channel
	signal rsp_xbar_demux_032_src0_ready                                                                : std_logic;                      -- rsp_xbar_mux_001:sink32_ready -> rsp_xbar_demux_032:src0_ready
	signal limiter_cmd_src_endofpacket                                                                  : std_logic;                      -- limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal limiter_cmd_src_startofpacket                                                                : std_logic;                      -- limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal limiter_cmd_src_data                                                                         : std_logic_vector(103 downto 0); -- limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	signal limiter_cmd_src_channel                                                                      : std_logic_vector(32 downto 0);  -- limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	signal limiter_cmd_src_ready                                                                        : std_logic;                      -- cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                 : std_logic;                      -- rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	signal rsp_xbar_mux_src_valid                                                                       : std_logic;                      -- rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	signal rsp_xbar_mux_src_startofpacket                                                               : std_logic;                      -- rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	signal rsp_xbar_mux_src_data                                                                        : std_logic_vector(103 downto 0); -- rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	signal rsp_xbar_mux_src_channel                                                                     : std_logic_vector(32 downto 0);  -- rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	signal rsp_xbar_mux_src_ready                                                                       : std_logic;                      -- limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	signal addr_router_001_src_endofpacket                                                              : std_logic;                      -- addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal addr_router_001_src_valid                                                                    : std_logic;                      -- addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	signal addr_router_001_src_startofpacket                                                            : std_logic;                      -- addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal addr_router_001_src_data                                                                     : std_logic_vector(103 downto 0); -- addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	signal addr_router_001_src_channel                                                                  : std_logic_vector(32 downto 0);  -- addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	signal addr_router_001_src_ready                                                                    : std_logic;                      -- cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                             : std_logic;                      -- rsp_xbar_mux_001:src_endofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                   : std_logic;                      -- rsp_xbar_mux_001:src_valid -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                           : std_logic;                      -- rsp_xbar_mux_001:src_startofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                    : std_logic_vector(103 downto 0); -- rsp_xbar_mux_001:src_data -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_001_src_channel                                                                 : std_logic_vector(32 downto 0);  -- rsp_xbar_mux_001:src_channel -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_001_src_ready                                                                   : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	signal cmd_xbar_mux_src_endofpacket                                                                 : std_logic;                      -- cmd_xbar_mux:src_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_src_valid                                                                       : std_logic;                      -- cmd_xbar_mux:src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_src_startofpacket                                                               : std_logic;                      -- cmd_xbar_mux:src_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_src_data                                                                        : std_logic_vector(103 downto 0); -- cmd_xbar_mux:src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_src_channel                                                                     : std_logic_vector(32 downto 0);  -- cmd_xbar_mux:src_channel -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_src_ready                                                                       : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                    : std_logic;                      -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                          : std_logic;                      -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                  : std_logic;                      -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                           : std_logic_vector(103 downto 0); -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                        : std_logic_vector(32 downto 0);  -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                          : std_logic;                      -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_mux_002_src_endofpacket                                                             : std_logic;                      -- cmd_xbar_mux_002:src_endofpacket -> system_id_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_002_src_valid                                                                   : std_logic;                      -- cmd_xbar_mux_002:src_valid -> system_id_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_002_src_startofpacket                                                           : std_logic;                      -- cmd_xbar_mux_002:src_startofpacket -> system_id_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_002_src_data                                                                    : std_logic_vector(103 downto 0); -- cmd_xbar_mux_002:src_data -> system_id_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_002_src_channel                                                                 : std_logic_vector(32 downto 0);  -- cmd_xbar_mux_002:src_channel -> system_id_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_002_src_ready                                                                   : std_logic;                      -- system_id_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	signal id_router_002_src_endofpacket                                                                : std_logic;                      -- id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal id_router_002_src_valid                                                                      : std_logic;                      -- id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	signal id_router_002_src_startofpacket                                                              : std_logic;                      -- id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal id_router_002_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	signal id_router_002_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	signal id_router_002_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	signal crosser_out_ready                                                                            : std_logic;                      -- pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	signal id_router_003_src_endofpacket                                                                : std_logic;                      -- id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal id_router_003_src_valid                                                                      : std_logic;                      -- id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	signal id_router_003_src_startofpacket                                                              : std_logic;                      -- id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal id_router_003_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	signal id_router_003_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	signal id_router_003_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	signal cmd_xbar_demux_001_src4_ready                                                                : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	signal id_router_004_src_endofpacket                                                                : std_logic;                      -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                      : std_logic;                      -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                              : std_logic;                      -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_demux_001_src5_ready                                                                : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	signal id_router_005_src_endofpacket                                                                : std_logic;                      -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                      : std_logic;                      -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                              : std_logic;                      -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal cmd_xbar_demux_001_src6_ready                                                                : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	signal id_router_006_src_endofpacket                                                                : std_logic;                      -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                      : std_logic;                      -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                              : std_logic;                      -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal cmd_xbar_demux_001_src7_ready                                                                : std_logic;                      -- pio_in_sw_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	signal id_router_007_src_endofpacket                                                                : std_logic;                      -- id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal id_router_007_src_valid                                                                      : std_logic;                      -- id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	signal id_router_007_src_startofpacket                                                              : std_logic;                      -- id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal id_router_007_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	signal id_router_007_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	signal id_router_007_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	signal cmd_xbar_demux_001_src8_ready                                                                : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	signal id_router_008_src_endofpacket                                                                : std_logic;                      -- id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	signal id_router_008_src_valid                                                                      : std_logic;                      -- id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	signal id_router_008_src_startofpacket                                                              : std_logic;                      -- id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	signal id_router_008_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	signal id_router_008_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	signal id_router_008_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	signal cmd_xbar_demux_001_src9_ready                                                                : std_logic;                      -- pio_in_ext_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	signal id_router_009_src_endofpacket                                                                : std_logic;                      -- id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	signal id_router_009_src_valid                                                                      : std_logic;                      -- id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	signal id_router_009_src_startofpacket                                                              : std_logic;                      -- id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	signal id_router_009_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	signal id_router_009_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	signal id_router_009_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	signal cmd_xbar_demux_001_src10_ready                                                               : std_logic;                      -- pio_out_red_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	signal id_router_010_src_endofpacket                                                                : std_logic;                      -- id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	signal id_router_010_src_valid                                                                      : std_logic;                      -- id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	signal id_router_010_src_startofpacket                                                              : std_logic;                      -- id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	signal id_router_010_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	signal id_router_010_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	signal id_router_010_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	signal cmd_xbar_demux_001_src11_ready                                                               : std_logic;                      -- pio_out_green_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	signal id_router_011_src_endofpacket                                                                : std_logic;                      -- id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	signal id_router_011_src_valid                                                                      : std_logic;                      -- id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	signal id_router_011_src_startofpacket                                                              : std_logic;                      -- id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	signal id_router_011_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	signal id_router_011_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	signal id_router_011_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	signal cmd_xbar_demux_001_src12_ready                                                               : std_logic;                      -- pio_out_ext_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	signal id_router_012_src_endofpacket                                                                : std_logic;                      -- id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	signal id_router_012_src_valid                                                                      : std_logic;                      -- id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	signal id_router_012_src_startofpacket                                                              : std_logic;                      -- id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	signal id_router_012_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	signal id_router_012_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	signal id_router_012_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	signal cmd_xbar_demux_001_src13_ready                                                               : std_logic;                      -- pio_async_reset_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	signal id_router_013_src_endofpacket                                                                : std_logic;                      -- id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	signal id_router_013_src_valid                                                                      : std_logic;                      -- id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	signal id_router_013_src_startofpacket                                                              : std_logic;                      -- id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	signal id_router_013_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	signal id_router_013_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	signal id_router_013_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	signal cmd_xbar_demux_001_src14_ready                                                               : std_logic;                      -- pio_en_mux_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src14_ready
	signal id_router_014_src_endofpacket                                                                : std_logic;                      -- id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	signal id_router_014_src_valid                                                                      : std_logic;                      -- id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	signal id_router_014_src_startofpacket                                                              : std_logic;                      -- id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	signal id_router_014_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	signal id_router_014_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	signal id_router_014_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	signal cmd_xbar_demux_001_src15_ready                                                               : std_logic;                      -- pio_direc_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src15_ready
	signal id_router_015_src_endofpacket                                                                : std_logic;                      -- id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	signal id_router_015_src_valid                                                                      : std_logic;                      -- id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	signal id_router_015_src_startofpacket                                                              : std_logic;                      -- id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	signal id_router_015_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	signal id_router_015_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	signal id_router_015_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	signal cmd_xbar_demux_001_src16_ready                                                               : std_logic;                      -- pio_direc_ram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src16_ready
	signal id_router_016_src_endofpacket                                                                : std_logic;                      -- id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	signal id_router_016_src_valid                                                                      : std_logic;                      -- id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	signal id_router_016_src_startofpacket                                                              : std_logic;                      -- id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	signal id_router_016_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	signal id_router_016_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	signal id_router_016_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	signal cmd_xbar_demux_001_src17_ready                                                               : std_logic;                      -- pio_wr_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src17_ready
	signal id_router_017_src_endofpacket                                                                : std_logic;                      -- id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	signal id_router_017_src_valid                                                                      : std_logic;                      -- id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	signal id_router_017_src_startofpacket                                                              : std_logic;                      -- id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	signal id_router_017_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	signal id_router_017_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	signal id_router_017_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	signal cmd_xbar_demux_001_src18_ready                                                               : std_logic;                      -- pio_sel_salida_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src18_ready
	signal id_router_018_src_endofpacket                                                                : std_logic;                      -- id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	signal id_router_018_src_valid                                                                      : std_logic;                      -- id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	signal id_router_018_src_startofpacket                                                              : std_logic;                      -- id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	signal id_router_018_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	signal id_router_018_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	signal id_router_018_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	signal cmd_xbar_demux_001_src19_ready                                                               : std_logic;                      -- pio_datos_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src19_ready
	signal id_router_019_src_endofpacket                                                                : std_logic;                      -- id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	signal id_router_019_src_valid                                                                      : std_logic;                      -- id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	signal id_router_019_src_startofpacket                                                              : std_logic;                      -- id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	signal id_router_019_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	signal id_router_019_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	signal id_router_019_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	signal cmd_xbar_demux_001_src20_ready                                                               : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src20_ready
	signal id_router_020_src_endofpacket                                                                : std_logic;                      -- id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	signal id_router_020_src_valid                                                                      : std_logic;                      -- id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	signal id_router_020_src_startofpacket                                                              : std_logic;                      -- id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	signal id_router_020_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	signal id_router_020_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	signal id_router_020_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	signal cmd_xbar_demux_001_src21_ready                                                               : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src21_ready
	signal id_router_021_src_endofpacket                                                                : std_logic;                      -- id_router_021:src_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	signal id_router_021_src_valid                                                                      : std_logic;                      -- id_router_021:src_valid -> rsp_xbar_demux_021:sink_valid
	signal id_router_021_src_startofpacket                                                              : std_logic;                      -- id_router_021:src_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	signal id_router_021_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_021:src_data -> rsp_xbar_demux_021:sink_data
	signal id_router_021_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_021:src_channel -> rsp_xbar_demux_021:sink_channel
	signal id_router_021_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_021:sink_ready -> id_router_021:src_ready
	signal cmd_xbar_demux_001_src22_ready                                                               : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src22_ready
	signal id_router_022_src_endofpacket                                                                : std_logic;                      -- id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	signal id_router_022_src_valid                                                                      : std_logic;                      -- id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	signal id_router_022_src_startofpacket                                                              : std_logic;                      -- id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	signal id_router_022_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	signal id_router_022_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	signal id_router_022_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	signal cmd_xbar_demux_001_src23_ready                                                               : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src23_ready
	signal id_router_023_src_endofpacket                                                                : std_logic;                      -- id_router_023:src_endofpacket -> rsp_xbar_demux_023:sink_endofpacket
	signal id_router_023_src_valid                                                                      : std_logic;                      -- id_router_023:src_valid -> rsp_xbar_demux_023:sink_valid
	signal id_router_023_src_startofpacket                                                              : std_logic;                      -- id_router_023:src_startofpacket -> rsp_xbar_demux_023:sink_startofpacket
	signal id_router_023_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_023:src_data -> rsp_xbar_demux_023:sink_data
	signal id_router_023_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_023:src_channel -> rsp_xbar_demux_023:sink_channel
	signal id_router_023_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_023:sink_ready -> id_router_023:src_ready
	signal cmd_xbar_demux_001_src24_ready                                                               : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src24_ready
	signal id_router_024_src_endofpacket                                                                : std_logic;                      -- id_router_024:src_endofpacket -> rsp_xbar_demux_024:sink_endofpacket
	signal id_router_024_src_valid                                                                      : std_logic;                      -- id_router_024:src_valid -> rsp_xbar_demux_024:sink_valid
	signal id_router_024_src_startofpacket                                                              : std_logic;                      -- id_router_024:src_startofpacket -> rsp_xbar_demux_024:sink_startofpacket
	signal id_router_024_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_024:src_data -> rsp_xbar_demux_024:sink_data
	signal id_router_024_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_024:src_channel -> rsp_xbar_demux_024:sink_channel
	signal id_router_024_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_024:sink_ready -> id_router_024:src_ready
	signal cmd_xbar_demux_001_src25_ready                                                               : std_logic;                      -- pio_captura_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src25_ready
	signal id_router_025_src_endofpacket                                                                : std_logic;                      -- id_router_025:src_endofpacket -> rsp_xbar_demux_025:sink_endofpacket
	signal id_router_025_src_valid                                                                      : std_logic;                      -- id_router_025:src_valid -> rsp_xbar_demux_025:sink_valid
	signal id_router_025_src_startofpacket                                                              : std_logic;                      -- id_router_025:src_startofpacket -> rsp_xbar_demux_025:sink_startofpacket
	signal id_router_025_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_025:src_data -> rsp_xbar_demux_025:sink_data
	signal id_router_025_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_025:src_channel -> rsp_xbar_demux_025:sink_channel
	signal id_router_025_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_025:sink_ready -> id_router_025:src_ready
	signal cmd_xbar_demux_001_src26_ready                                                               : std_logic;                      -- pio_captura_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src26_ready
	signal id_router_026_src_endofpacket                                                                : std_logic;                      -- id_router_026:src_endofpacket -> rsp_xbar_demux_026:sink_endofpacket
	signal id_router_026_src_valid                                                                      : std_logic;                      -- id_router_026:src_valid -> rsp_xbar_demux_026:sink_valid
	signal id_router_026_src_startofpacket                                                              : std_logic;                      -- id_router_026:src_startofpacket -> rsp_xbar_demux_026:sink_startofpacket
	signal id_router_026_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_026:src_data -> rsp_xbar_demux_026:sink_data
	signal id_router_026_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_026:src_channel -> rsp_xbar_demux_026:sink_channel
	signal id_router_026_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_026:sink_ready -> id_router_026:src_ready
	signal cmd_xbar_demux_001_src27_ready                                                               : std_logic;                      -- pio_captura_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src27_ready
	signal id_router_027_src_endofpacket                                                                : std_logic;                      -- id_router_027:src_endofpacket -> rsp_xbar_demux_027:sink_endofpacket
	signal id_router_027_src_valid                                                                      : std_logic;                      -- id_router_027:src_valid -> rsp_xbar_demux_027:sink_valid
	signal id_router_027_src_startofpacket                                                              : std_logic;                      -- id_router_027:src_startofpacket -> rsp_xbar_demux_027:sink_startofpacket
	signal id_router_027_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_027:src_data -> rsp_xbar_demux_027:sink_data
	signal id_router_027_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_027:src_channel -> rsp_xbar_demux_027:sink_channel
	signal id_router_027_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_027:sink_ready -> id_router_027:src_ready
	signal cmd_xbar_demux_001_src28_ready                                                               : std_logic;                      -- pio_captura_3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src28_ready
	signal id_router_028_src_endofpacket                                                                : std_logic;                      -- id_router_028:src_endofpacket -> rsp_xbar_demux_028:sink_endofpacket
	signal id_router_028_src_valid                                                                      : std_logic;                      -- id_router_028:src_valid -> rsp_xbar_demux_028:sink_valid
	signal id_router_028_src_startofpacket                                                              : std_logic;                      -- id_router_028:src_startofpacket -> rsp_xbar_demux_028:sink_startofpacket
	signal id_router_028_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_028:src_data -> rsp_xbar_demux_028:sink_data
	signal id_router_028_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_028:src_channel -> rsp_xbar_demux_028:sink_channel
	signal id_router_028_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_028:sink_ready -> id_router_028:src_ready
	signal cmd_xbar_demux_001_src29_ready                                                               : std_logic;                      -- pio_captura_4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src29_ready
	signal id_router_029_src_endofpacket                                                                : std_logic;                      -- id_router_029:src_endofpacket -> rsp_xbar_demux_029:sink_endofpacket
	signal id_router_029_src_valid                                                                      : std_logic;                      -- id_router_029:src_valid -> rsp_xbar_demux_029:sink_valid
	signal id_router_029_src_startofpacket                                                              : std_logic;                      -- id_router_029:src_startofpacket -> rsp_xbar_demux_029:sink_startofpacket
	signal id_router_029_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_029:src_data -> rsp_xbar_demux_029:sink_data
	signal id_router_029_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_029:src_channel -> rsp_xbar_demux_029:sink_channel
	signal id_router_029_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_029:sink_ready -> id_router_029:src_ready
	signal cmd_xbar_demux_001_src30_ready                                                               : std_logic;                      -- pio_in_32_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src30_ready
	signal id_router_030_src_endofpacket                                                                : std_logic;                      -- id_router_030:src_endofpacket -> rsp_xbar_demux_030:sink_endofpacket
	signal id_router_030_src_valid                                                                      : std_logic;                      -- id_router_030:src_valid -> rsp_xbar_demux_030:sink_valid
	signal id_router_030_src_startofpacket                                                              : std_logic;                      -- id_router_030:src_startofpacket -> rsp_xbar_demux_030:sink_startofpacket
	signal id_router_030_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_030:src_data -> rsp_xbar_demux_030:sink_data
	signal id_router_030_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_030:src_channel -> rsp_xbar_demux_030:sink_channel
	signal id_router_030_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_030:sink_ready -> id_router_030:src_ready
	signal cmd_xbar_demux_001_src31_ready                                                               : std_logic;                      -- lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src31_ready
	signal id_router_031_src_endofpacket                                                                : std_logic;                      -- id_router_031:src_endofpacket -> rsp_xbar_demux_031:sink_endofpacket
	signal id_router_031_src_valid                                                                      : std_logic;                      -- id_router_031:src_valid -> rsp_xbar_demux_031:sink_valid
	signal id_router_031_src_startofpacket                                                              : std_logic;                      -- id_router_031:src_startofpacket -> rsp_xbar_demux_031:sink_startofpacket
	signal id_router_031_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_031:src_data -> rsp_xbar_demux_031:sink_data
	signal id_router_031_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_031:src_channel -> rsp_xbar_demux_031:sink_channel
	signal id_router_031_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_031:sink_ready -> id_router_031:src_ready
	signal cmd_xbar_demux_001_src32_ready                                                               : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src32_ready
	signal id_router_032_src_endofpacket                                                                : std_logic;                      -- id_router_032:src_endofpacket -> rsp_xbar_demux_032:sink_endofpacket
	signal id_router_032_src_valid                                                                      : std_logic;                      -- id_router_032:src_valid -> rsp_xbar_demux_032:sink_valid
	signal id_router_032_src_startofpacket                                                              : std_logic;                      -- id_router_032:src_startofpacket -> rsp_xbar_demux_032:sink_startofpacket
	signal id_router_032_src_data                                                                       : std_logic_vector(103 downto 0); -- id_router_032:src_data -> rsp_xbar_demux_032:sink_data
	signal id_router_032_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_032:src_channel -> rsp_xbar_demux_032:sink_channel
	signal id_router_032_src_ready                                                                      : std_logic;                      -- rsp_xbar_demux_032:sink_ready -> id_router_032:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                             : std_logic;                      -- cmd_xbar_mux_001:src_endofpacket -> width_adapter:in_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                   : std_logic;                      -- cmd_xbar_mux_001:src_valid -> width_adapter:in_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                           : std_logic;                      -- cmd_xbar_mux_001:src_startofpacket -> width_adapter:in_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                    : std_logic_vector(103 downto 0); -- cmd_xbar_mux_001:src_data -> width_adapter:in_data
	signal cmd_xbar_mux_001_src_channel                                                                 : std_logic_vector(32 downto 0);  -- cmd_xbar_mux_001:src_channel -> width_adapter:in_channel
	signal cmd_xbar_mux_001_src_ready                                                                   : std_logic;                      -- width_adapter:in_ready -> cmd_xbar_mux_001:src_ready
	signal width_adapter_src_endofpacket                                                                : std_logic;                      -- width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	signal width_adapter_src_valid                                                                      : std_logic;                      -- width_adapter:out_valid -> burst_adapter:sink0_valid
	signal width_adapter_src_startofpacket                                                              : std_logic;                      -- width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	signal width_adapter_src_data                                                                       : std_logic_vector(85 downto 0);  -- width_adapter:out_data -> burst_adapter:sink0_data
	signal width_adapter_src_ready                                                                      : std_logic;                      -- burst_adapter:sink0_ready -> width_adapter:out_ready
	signal width_adapter_src_channel                                                                    : std_logic_vector(32 downto 0);  -- width_adapter:out_channel -> burst_adapter:sink0_channel
	signal id_router_001_src_endofpacket                                                                : std_logic;                      -- id_router_001:src_endofpacket -> width_adapter_001:in_endofpacket
	signal id_router_001_src_valid                                                                      : std_logic;                      -- id_router_001:src_valid -> width_adapter_001:in_valid
	signal id_router_001_src_startofpacket                                                              : std_logic;                      -- id_router_001:src_startofpacket -> width_adapter_001:in_startofpacket
	signal id_router_001_src_data                                                                       : std_logic_vector(85 downto 0);  -- id_router_001:src_data -> width_adapter_001:in_data
	signal id_router_001_src_channel                                                                    : std_logic_vector(32 downto 0);  -- id_router_001:src_channel -> width_adapter_001:in_channel
	signal id_router_001_src_ready                                                                      : std_logic;                      -- width_adapter_001:in_ready -> id_router_001:src_ready
	signal width_adapter_001_src_endofpacket                                                            : std_logic;                      -- width_adapter_001:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal width_adapter_001_src_valid                                                                  : std_logic;                      -- width_adapter_001:out_valid -> rsp_xbar_demux_001:sink_valid
	signal width_adapter_001_src_startofpacket                                                          : std_logic;                      -- width_adapter_001:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal width_adapter_001_src_data                                                                   : std_logic_vector(103 downto 0); -- width_adapter_001:out_data -> rsp_xbar_demux_001:sink_data
	signal width_adapter_001_src_ready                                                                  : std_logic;                      -- rsp_xbar_demux_001:sink_ready -> width_adapter_001:out_ready
	signal width_adapter_001_src_channel                                                                : std_logic_vector(32 downto 0);  -- width_adapter_001:out_channel -> rsp_xbar_demux_001:sink_channel
	signal crosser_out_endofpacket                                                                      : std_logic;                      -- crosser:out_endofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal crosser_out_valid                                                                            : std_logic;                      -- crosser:out_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal crosser_out_startofpacket                                                                    : std_logic;                      -- crosser:out_startofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal crosser_out_data                                                                             : std_logic_vector(103 downto 0); -- crosser:out_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal crosser_out_channel                                                                          : std_logic_vector(32 downto 0);  -- crosser:out_channel -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src3_endofpacket                                                          : std_logic;                      -- cmd_xbar_demux_001:src3_endofpacket -> crosser:in_endofpacket
	signal cmd_xbar_demux_001_src3_valid                                                                : std_logic;                      -- cmd_xbar_demux_001:src3_valid -> crosser:in_valid
	signal cmd_xbar_demux_001_src3_startofpacket                                                        : std_logic;                      -- cmd_xbar_demux_001:src3_startofpacket -> crosser:in_startofpacket
	signal cmd_xbar_demux_001_src3_data                                                                 : std_logic_vector(103 downto 0); -- cmd_xbar_demux_001:src3_data -> crosser:in_data
	signal cmd_xbar_demux_001_src3_channel                                                              : std_logic_vector(32 downto 0);  -- cmd_xbar_demux_001:src3_channel -> crosser:in_channel
	signal cmd_xbar_demux_001_src3_ready                                                                : std_logic;                      -- crosser:in_ready -> cmd_xbar_demux_001:src3_ready
	signal crosser_001_out_endofpacket                                                                  : std_logic;                      -- crosser_001:out_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	signal crosser_001_out_valid                                                                        : std_logic;                      -- crosser_001:out_valid -> rsp_xbar_mux_001:sink3_valid
	signal crosser_001_out_startofpacket                                                                : std_logic;                      -- crosser_001:out_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	signal crosser_001_out_data                                                                         : std_logic_vector(103 downto 0); -- crosser_001:out_data -> rsp_xbar_mux_001:sink3_data
	signal crosser_001_out_channel                                                                      : std_logic_vector(32 downto 0);  -- crosser_001:out_channel -> rsp_xbar_mux_001:sink3_channel
	signal crosser_001_out_ready                                                                        : std_logic;                      -- rsp_xbar_mux_001:sink3_ready -> crosser_001:out_ready
	signal rsp_xbar_demux_003_src0_endofpacket                                                          : std_logic;                      -- rsp_xbar_demux_003:src0_endofpacket -> crosser_001:in_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                : std_logic;                      -- rsp_xbar_demux_003:src0_valid -> crosser_001:in_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                        : std_logic;                      -- rsp_xbar_demux_003:src0_startofpacket -> crosser_001:in_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                 : std_logic_vector(103 downto 0); -- rsp_xbar_demux_003:src0_data -> crosser_001:in_data
	signal rsp_xbar_demux_003_src0_channel                                                              : std_logic_vector(32 downto 0);  -- rsp_xbar_demux_003:src0_channel -> crosser_001:in_channel
	signal rsp_xbar_demux_003_src0_ready                                                                : std_logic;                      -- crosser_001:in_ready -> rsp_xbar_demux_003:src0_ready
	signal limiter_cmd_valid_data                                                                       : std_logic_vector(32 downto 0);  -- limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	signal irq_mapper_receiver0_irq                                                                     : std_logic;                      -- pio_captura_3:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                                     : std_logic;                      -- pio_captura_2:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                                     : std_logic;                      -- pio_in_ext:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                                                     : std_logic;                      -- uart:av_irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                                                     : std_logic;                      -- timer_0:irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                                                     : std_logic;                      -- timer_1:irq -> irq_mapper:receiver5_irq
	signal irq_mapper_receiver6_irq                                                                     : std_logic;                      -- pio_in_key_edge:irq -> irq_mapper:receiver6_irq
	signal irq_mapper_receiver7_irq                                                                     : std_logic;                      -- pio_compara_int_0:irq -> irq_mapper:receiver7_irq
	signal irq_mapper_receiver8_irq                                                                     : std_logic;                      -- pio_compara_int_1:irq -> irq_mapper:receiver8_irq
	signal irq_mapper_receiver9_irq                                                                     : std_logic;                      -- pio_compara_int_2:irq -> irq_mapper:receiver9_irq
	signal irq_mapper_receiver10_irq                                                                    : std_logic;                      -- pio_compara_int_3:irq -> irq_mapper:receiver10_irq
	signal irq_mapper_receiver11_irq                                                                    : std_logic;                      -- pio_compara_int_4:irq -> irq_mapper:receiver11_irq
	signal irq_mapper_receiver12_irq                                                                    : std_logic;                      -- pio_captura_0:irq -> irq_mapper:receiver12_irq
	signal irq_mapper_receiver13_irq                                                                    : std_logic;                      -- pio_captura_1:irq -> irq_mapper:receiver13_irq
	signal irq_mapper_receiver14_irq                                                                    : std_logic;                      -- pio_captura_4:irq -> irq_mapper:receiver14_irq
	signal irq_mapper_receiver15_irq                                                                    : std_logic;                      -- DM9000A:oINT -> irq_mapper:receiver15_irq
	signal cpu_d_irq_irq                                                                                : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> cpu:d_irq
	signal reset_reset_n_ports_inv                                                                      : std_logic;                      -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal sdram_s1_translator_avalon_anti_slave_0_write_ports_inv                                      : std_logic;                      -- sdram_s1_translator_avalon_anti_slave_0_write:inv -> sdram:az_wr_n
	signal sdram_s1_translator_avalon_anti_slave_0_read_ports_inv                                       : std_logic;                      -- sdram_s1_translator_avalon_anti_slave_0_read:inv -> sdram:az_rd_n
	signal sdram_s1_translator_avalon_anti_slave_0_byteenable_ports_inv                                 : std_logic_vector(1 downto 0);   -- sdram_s1_translator_avalon_anti_slave_0_byteenable:inv -> sdram:az_be_n
	signal uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                        : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> uart:av_write_n
	signal uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                         : std_logic;                      -- uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> uart:av_read_n
	signal timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv                                    : std_logic;                      -- timer_0_s1_translator_avalon_anti_slave_0_write:inv -> timer_0:write_n
	signal timer_1_s1_translator_avalon_anti_slave_0_write_ports_inv                                    : std_logic;                      -- timer_1_s1_translator_avalon_anti_slave_0_write:inv -> timer_1:write_n
	signal pio_in_key_edge_s1_translator_avalon_anti_slave_0_write_ports_inv                            : std_logic;                      -- pio_in_key_edge_s1_translator_avalon_anti_slave_0_write:inv -> pio_in_key_edge:write_n
	signal pio_in_ext_s1_translator_avalon_anti_slave_0_write_ports_inv                                 : std_logic;                      -- pio_in_ext_s1_translator_avalon_anti_slave_0_write:inv -> pio_in_ext:write_n
	signal pio_out_red_s1_translator_avalon_anti_slave_0_write_ports_inv                                : std_logic;                      -- pio_out_red_s1_translator_avalon_anti_slave_0_write:inv -> pio_out_red:write_n
	signal pio_out_green_s1_translator_avalon_anti_slave_0_write_ports_inv                              : std_logic;                      -- pio_out_green_s1_translator_avalon_anti_slave_0_write:inv -> pio_out_green:write_n
	signal pio_out_ext_s1_translator_avalon_anti_slave_0_write_ports_inv                                : std_logic;                      -- pio_out_ext_s1_translator_avalon_anti_slave_0_write:inv -> pio_out_ext:write_n
	signal pio_async_reset_s1_translator_avalon_anti_slave_0_write_ports_inv                            : std_logic;                      -- pio_async_reset_s1_translator_avalon_anti_slave_0_write:inv -> pio_async_reset:write_n
	signal pio_en_mux_s1_translator_avalon_anti_slave_0_write_ports_inv                                 : std_logic;                      -- pio_en_mux_s1_translator_avalon_anti_slave_0_write:inv -> pio_en_mux:write_n
	signal pio_direc_s1_translator_avalon_anti_slave_0_write_ports_inv                                  : std_logic;                      -- pio_direc_s1_translator_avalon_anti_slave_0_write:inv -> pio_direc:write_n
	signal pio_direc_ram_s1_translator_avalon_anti_slave_0_write_ports_inv                              : std_logic;                      -- pio_direc_ram_s1_translator_avalon_anti_slave_0_write:inv -> pio_direc_ram:write_n
	signal pio_wr_s1_translator_avalon_anti_slave_0_write_ports_inv                                     : std_logic;                      -- pio_wr_s1_translator_avalon_anti_slave_0_write:inv -> pio_wr:write_n
	signal pio_sel_salida_s1_translator_avalon_anti_slave_0_write_ports_inv                             : std_logic;                      -- pio_sel_salida_s1_translator_avalon_anti_slave_0_write:inv -> pio_sel_salida:write_n
	signal pio_datos_s1_translator_avalon_anti_slave_0_write_ports_inv                                  : std_logic;                      -- pio_datos_s1_translator_avalon_anti_slave_0_write:inv -> pio_datos:write_n
	signal pio_compara_int_0_s1_translator_avalon_anti_slave_0_write_ports_inv                          : std_logic;                      -- pio_compara_int_0_s1_translator_avalon_anti_slave_0_write:inv -> pio_compara_int_0:write_n
	signal pio_compara_int_1_s1_translator_avalon_anti_slave_0_write_ports_inv                          : std_logic;                      -- pio_compara_int_1_s1_translator_avalon_anti_slave_0_write:inv -> pio_compara_int_1:write_n
	signal pio_compara_int_2_s1_translator_avalon_anti_slave_0_write_ports_inv                          : std_logic;                      -- pio_compara_int_2_s1_translator_avalon_anti_slave_0_write:inv -> pio_compara_int_2:write_n
	signal pio_compara_int_3_s1_translator_avalon_anti_slave_0_write_ports_inv                          : std_logic;                      -- pio_compara_int_3_s1_translator_avalon_anti_slave_0_write:inv -> pio_compara_int_3:write_n
	signal pio_compara_int_4_s1_translator_avalon_anti_slave_0_write_ports_inv                          : std_logic;                      -- pio_compara_int_4_s1_translator_avalon_anti_slave_0_write:inv -> pio_compara_int_4:write_n
	signal pio_captura_0_s1_translator_avalon_anti_slave_0_write_ports_inv                              : std_logic;                      -- pio_captura_0_s1_translator_avalon_anti_slave_0_write:inv -> pio_captura_0:write_n
	signal pio_captura_1_s1_translator_avalon_anti_slave_0_write_ports_inv                              : std_logic;                      -- pio_captura_1_s1_translator_avalon_anti_slave_0_write:inv -> pio_captura_1:write_n
	signal pio_captura_2_s1_translator_avalon_anti_slave_0_write_ports_inv                              : std_logic;                      -- pio_captura_2_s1_translator_avalon_anti_slave_0_write:inv -> pio_captura_2:write_n
	signal pio_captura_3_s1_translator_avalon_anti_slave_0_write_ports_inv                              : std_logic;                      -- pio_captura_3_s1_translator_avalon_anti_slave_0_write:inv -> pio_captura_3:write_n
	signal pio_captura_4_s1_translator_avalon_anti_slave_0_write_ports_inv                              : std_logic;                      -- pio_captura_4_s1_translator_avalon_anti_slave_0_write:inv -> pio_captura_4:write_n
	signal pio_in_32_s1_translator_avalon_anti_slave_0_write_ports_inv                                  : std_logic;                      -- pio_in_32_s1_translator_avalon_anti_slave_0_write:inv -> pio_in_32:write_n
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect_ports_inv                   : std_logic;                      -- dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect:inv -> DM9000A:iCS_N
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write_ports_inv                        : std_logic;                      -- dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write:inv -> DM9000A:iWR_N
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read_ports_inv                         : std_logic;                      -- dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read:inv -> DM9000A:iRD_N
	signal rst_controller_reset_out_reset_ports_inv                                                     : std_logic;                      -- rst_controller_reset_out_reset:inv -> [DM9000A:iRST_N, cpu:reset_n, lcd:reset_n, pio_async_reset:reset_n, pio_captura_0:reset_n, pio_captura_1:reset_n, pio_captura_2:reset_n, pio_captura_3:reset_n, pio_captura_4:reset_n, pio_compara_int_0:reset_n, pio_compara_int_1:reset_n, pio_compara_int_2:reset_n, pio_compara_int_3:reset_n, pio_compara_int_4:reset_n, pio_datos:reset_n, pio_direc:reset_n, pio_direc_ram:reset_n, pio_en_mux:reset_n, pio_in_32:reset_n, pio_in_ext:reset_n, pio_in_key_edge:reset_n, pio_in_sw:reset_n, pio_out_ext:reset_n, pio_out_green:reset_n, pio_out_red:reset_n, pio_sel_salida:reset_n, pio_wr:reset_n, sdram:reset_n, system_id:reset_n, timer_0:reset_n, timer_1:reset_n, uart:rst_n]

begin

	cpu : component NIOSIImicro_cpu
		port map (
			clk                                   => pll_c0_clk,                                                       --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                         --                   reset_n.reset_n
			d_address                             => cpu_data_master_address,                                          --               data_master.address
			d_byteenable                          => cpu_data_master_byteenable,                                       --                          .byteenable
			d_read                                => cpu_data_master_read,                                             --                          .read
			d_readdata                            => cpu_data_master_readdata,                                         --                          .readdata
			d_waitrequest                         => cpu_data_master_waitrequest,                                      --                          .waitrequest
			d_write                               => cpu_data_master_write,                                            --                          .write
			d_writedata                           => cpu_data_master_writedata,                                        --                          .writedata
			jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,                                      --                          .debugaccess
			i_address                             => cpu_instruction_master_address,                                   --        instruction_master.address
			i_read                                => cpu_instruction_master_read,                                      --                          .read
			i_readdata                            => cpu_instruction_master_readdata,                                  --                          .readdata
			i_waitrequest                         => cpu_instruction_master_waitrequest,                               --                          .waitrequest
			i_readdatavalid                       => cpu_instruction_master_readdatavalid,                             --                          .readdatavalid
			d_irq                                 => cpu_d_irq_irq,                                                    --                     d_irq.irq
			jtag_debug_module_resetrequest        => open,                                                             --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => cpu_jtag_debug_module_translator_avalon_anti_slave_0_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => cpu_jtag_debug_module_translator_avalon_anti_slave_0_read,        --                          .read
			jtag_debug_module_readdata            => cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => cpu_jtag_debug_module_translator_avalon_anti_slave_0_write,       --                          .write
			jtag_debug_module_writedata           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata,   --                          .writedata
			no_ci_readra                          => open                                                              -- custom_instruction_master.readra
		);

	pll : component NIOSIImicro_pll
		port map (
			clk       => clk_50_clk,                                             --       inclk_interface.clk
			reset     => rst_controller_001_reset_out_reset,                     -- inclk_interface_reset.reset
			read      => pll_pll_slave_translator_avalon_anti_slave_0_read,      --             pll_slave.read
			write     => pll_pll_slave_translator_avalon_anti_slave_0_write,     --                      .write
			address   => pll_pll_slave_translator_avalon_anti_slave_0_address,   --                      .address
			readdata  => pll_pll_slave_translator_avalon_anti_slave_0_readdata,  --                      .readdata
			writedata => pll_pll_slave_translator_avalon_anti_slave_0_writedata, --                      .writedata
			c0        => pll_c0_clk,                                             --                    c0.clk
			c1        => clock_100_clk,                                          --                    c1.clk
			c2        => sdram_clock_clk,                                        --                    c2.clk
			areset    => open,                                                   --        areset_conduit.export
			locked    => open,                                                   --        locked_conduit.export
			phasedone => open                                                    --     phasedone_conduit.export
		);

	sdram : component NIOSIImicro_sdram
		port map (
			clk            => pll_c0_clk,                                                   --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                     -- reset.reset_n
			az_addr        => sdram_s1_translator_avalon_anti_slave_0_address,              --    s1.address
			az_be_n        => sdram_s1_translator_avalon_anti_slave_0_byteenable_ports_inv, --      .byteenable_n
			az_cs          => sdram_s1_translator_avalon_anti_slave_0_chipselect,           --      .chipselect
			az_data        => sdram_s1_translator_avalon_anti_slave_0_writedata,            --      .writedata
			az_rd_n        => sdram_s1_translator_avalon_anti_slave_0_read_ports_inv,       --      .read_n
			az_wr_n        => sdram_s1_translator_avalon_anti_slave_0_write_ports_inv,      --      .write_n
			za_data        => sdram_s1_translator_avalon_anti_slave_0_readdata,             --      .readdata
			za_valid       => sdram_s1_translator_avalon_anti_slave_0_readdatavalid,        --      .readdatavalid
			za_waitrequest => sdram_s1_translator_avalon_anti_slave_0_waitrequest,          --      .waitrequest
			zs_addr        => sdram_controller_addr,                                        --  wire.export
			zs_ba          => sdram_controller_ba,                                          --      .export
			zs_cas_n       => sdram_controller_cas_n,                                       --      .export
			zs_cke         => sdram_controller_cke,                                         --      .export
			zs_cs_n        => sdram_controller_cs_n,                                        --      .export
			zs_dq          => sdram_controller_dq,                                          --      .export
			zs_dqm         => sdram_controller_dqm,                                         --      .export
			zs_ras_n       => sdram_controller_ras_n,                                       --      .export
			zs_we_n        => sdram_controller_we_n                                         --      .export
		);

	uart : component NIOSIImicro_uart
		port map (
			clk            => pll_c0_clk,                                                            --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                              --             reset.reset_n
			av_chipselect  => uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address(0),      --                  .address
			av_read_n      => uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver3_irq                                               --               irq.irq
		);

	timer_0 : component NIOSIImicro_timer_0
		port map (
			clk        => pll_c0_clk,                                                --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  -- reset.reset_n
			address    => timer_0_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => timer_0_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => timer_0_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => timer_0_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver4_irq                                   --   irq.irq
		);

	timer_1 : component NIOSIImicro_timer_1
		port map (
			clk        => pll_c0_clk,                                                --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  -- reset.reset_n
			address    => timer_1_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => timer_1_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => timer_1_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => timer_1_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => timer_1_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver5_irq                                   --   irq.irq
		);

	pio_in_sw : component NIOSIImicro_pio_in_sw
		port map (
			clk      => pll_c0_clk,                                           --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,             --               reset.reset_n
			address  => pio_in_sw_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => pio_in_sw_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => pio_in_sw_export                                      -- external_connection.export
		);

	pio_in_key_edge : component NIOSIImicro_pio_in_key_edge
		port map (
			clk        => pll_c0_clk,                                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                          --               reset.reset_n
			address    => pio_in_key_edge_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_in_key_edge_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_in_key_edge_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_in_key_edge_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_in_key_edge_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => pio_in_key_edge_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver6_irq                                           --                 irq.irq
		);

	pio_in_ext : component NIOSIImicro_pio_in_ext
		port map (
			clk        => pll_c0_clk,                                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                     --               reset.reset_n
			address    => pio_in_ext_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_in_ext_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_in_ext_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_in_ext_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_in_ext_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => pio_in_ext_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver2_irq                                      --                 irq.irq
		);

	pio_out_red : component NIOSIImicro_pio_out_red
		port map (
			clk        => pll_c0_clk,                                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                      --               reset.reset_n
			address    => pio_out_red_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_out_red_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_out_red_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_out_red_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_out_red_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pio_out_red_export                                             -- external_connection.export
		);

	pio_out_green : component NIOSIImicro_pio_out_green
		port map (
			clk        => pll_c0_clk,                                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                        --               reset.reset_n
			address    => pio_out_green_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_out_green_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_out_green_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_out_green_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_out_green_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pio_out_green_export                                             -- external_connection.export
		);

	pio_out_ext : component NIOSIImicro_pio_out_ext
		port map (
			clk        => pll_c0_clk,                                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                      --               reset.reset_n
			address    => pio_out_ext_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_out_ext_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_out_ext_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_out_ext_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_out_ext_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pio_out_ext_export                                             -- external_connection.export
		);

	pio_en_mux : component NIOSIImicro_pio_en_mux
		port map (
			clk        => pll_c0_clk,                                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                     --               reset.reset_n
			address    => pio_en_mux_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_en_mux_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_en_mux_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_en_mux_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_en_mux_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pio_en_mux_export                                             -- external_connection.export
		);

	pio_direc : component NIOSIImicro_pio_direc
		port map (
			clk        => pll_c0_clk,                                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                    --               reset.reset_n
			address    => pio_direc_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_direc_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_direc_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_direc_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_direc_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pio_direc_export                                             -- external_connection.export
		);

	pio_direc_ram : component NIOSIImicro_pio_direc_ram
		port map (
			clk        => pll_c0_clk,                                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                        --               reset.reset_n
			address    => pio_direc_ram_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_direc_ram_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_direc_ram_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_direc_ram_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_direc_ram_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pio_direc_ram_export                                             -- external_connection.export
		);

	pio_wr : component NIOSIImicro_pio_en_mux
		port map (
			clk        => pll_c0_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                 --               reset.reset_n
			address    => pio_wr_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_wr_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_wr_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_wr_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_wr_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pio_wr_export                                             -- external_connection.export
		);

	pio_sel_salida : component NIOSIImicro_pio_direc
		port map (
			clk        => pll_c0_clk,                                                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                         --               reset.reset_n
			address    => pio_sel_salida_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_sel_salida_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_sel_salida_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_sel_salida_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_sel_salida_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pio_sel_salida_export                                             -- external_connection.export
		);

	pio_datos : component NIOSIImicro_pio_datos
		port map (
			clk        => pll_c0_clk,                                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                    --               reset.reset_n
			address    => pio_datos_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_datos_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_datos_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_datos_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_datos_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pio_datos_export                                             -- external_connection.export
		);

	pio_compara_int_0 : component NIOSIImicro_pio_compara_int_0
		port map (
			clk        => pll_c0_clk,                                                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                            --               reset.reset_n
			address    => pio_compara_int_0_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_compara_int_0_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_compara_int_0_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_compara_int_0_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_compara_int_0_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => pio_compara_int_0_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver7_irq                                             --                 irq.irq
		);

	pio_compara_int_1 : component NIOSIImicro_pio_compara_int_0
		port map (
			clk        => pll_c0_clk,                                                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                            --               reset.reset_n
			address    => pio_compara_int_1_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_compara_int_1_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_compara_int_1_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_compara_int_1_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_compara_int_1_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => pio_compara_int_1_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver8_irq                                             --                 irq.irq
		);

	pio_compara_int_2 : component NIOSIImicro_pio_compara_int_0
		port map (
			clk        => pll_c0_clk,                                                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                            --               reset.reset_n
			address    => pio_compara_int_2_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_compara_int_2_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_compara_int_2_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_compara_int_2_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_compara_int_2_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => pio_compara_int_2_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver9_irq                                             --                 irq.irq
		);

	pio_compara_int_3 : component NIOSIImicro_pio_compara_int_0
		port map (
			clk        => pll_c0_clk,                                                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                            --               reset.reset_n
			address    => pio_compara_int_3_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_compara_int_3_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_compara_int_3_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_compara_int_3_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_compara_int_3_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => pio_compara_int_3_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver10_irq                                            --                 irq.irq
		);

	pio_compara_int_4 : component NIOSIImicro_pio_compara_int_0
		port map (
			clk        => pll_c0_clk,                                                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                            --               reset.reset_n
			address    => pio_compara_int_4_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_compara_int_4_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_compara_int_4_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_compara_int_4_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_compara_int_4_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => pio_compara_int_4_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver11_irq                                            --                 irq.irq
		);

	pio_captura_0 : component NIOSIImicro_pio_compara_int_0
		port map (
			clk        => pll_c0_clk,                                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                        --               reset.reset_n
			address    => pio_captura_0_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_captura_0_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_captura_0_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_captura_0_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_captura_0_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => pio_captura_0_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver12_irq                                        --                 irq.irq
		);

	pio_captura_1 : component NIOSIImicro_pio_compara_int_0
		port map (
			clk        => pll_c0_clk,                                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                        --               reset.reset_n
			address    => pio_captura_1_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_captura_1_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_captura_1_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_captura_1_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_captura_1_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => pio_captura_1_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver13_irq                                        --                 irq.irq
		);

	pio_captura_2 : component NIOSIImicro_pio_compara_int_0
		port map (
			clk        => pll_c0_clk,                                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                        --               reset.reset_n
			address    => pio_captura_2_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_captura_2_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_captura_2_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_captura_2_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_captura_2_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => pio_captura_2_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver1_irq                                         --                 irq.irq
		);

	pio_captura_3 : component NIOSIImicro_pio_compara_int_0
		port map (
			clk        => pll_c0_clk,                                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                        --               reset.reset_n
			address    => pio_captura_3_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_captura_3_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_captura_3_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_captura_3_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_captura_3_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => pio_captura_3_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver0_irq                                         --                 irq.irq
		);

	pio_captura_4 : component NIOSIImicro_pio_compara_int_0
		port map (
			clk        => pll_c0_clk,                                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                        --               reset.reset_n
			address    => pio_captura_4_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_captura_4_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_captura_4_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_captura_4_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_captura_4_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => pio_captura_4_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver14_irq                                        --                 irq.irq
		);

	pio_in_32 : component NIOSIImicro_pio_in_32
		port map (
			clk        => pll_c0_clk,                                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                    --               reset.reset_n
			address    => pio_in_32_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_in_32_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_in_32_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_in_32_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_in_32_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => pio_in_32_export                                             -- external_connection.export
		);

	lcd : component NIOSIImicro_lcd
		port map (
			reset_n       => rst_controller_reset_out_reset_ports_inv,                       --         reset.reset_n
			clk           => pll_c0_clk,                                                     --           clk.clk
			begintransfer => lcd_control_slave_translator_avalon_anti_slave_0_begintransfer, -- control_slave.begintransfer
			read          => lcd_control_slave_translator_avalon_anti_slave_0_read,          --              .read
			write         => lcd_control_slave_translator_avalon_anti_slave_0_write,         --              .write
			readdata      => lcd_control_slave_translator_avalon_anti_slave_0_readdata,      --              .readdata
			writedata     => lcd_control_slave_translator_avalon_anti_slave_0_writedata,     --              .writedata
			address       => lcd_control_slave_translator_avalon_anti_slave_0_address,       --              .address
			LCD_RS        => lcd_RS,                                                         --      external.export
			LCD_RW        => lcd_RW,                                                         --              .export
			LCD_data      => lcd_data,                                                       --              .export
			LCD_E         => lcd_E                                                           --              .export
		);

	system_id : component NIOSIImicro_system_id
		port map (
			clock    => pll_c0_clk,                                                        --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                          --         reset.reset_n
			readdata => system_id_control_slave_translator_avalon_anti_slave_0_readdata,   -- control_slave.readdata
			address  => system_id_control_slave_translator_avalon_anti_slave_0_address(0)  --              .address
		);

	dm9000a : component DM9000A_IF
		port map (
			iCLK       => pll_c0_clk,                                                                 --                   clk.clk
			iRST_N     => rst_controller_reset_out_reset_ports_inv,                                   --             clk_reset.reset_n
			iOSC_50    => dm9000a_iOSC_50,                                                            -- avalon_slave_0_export.export
			ENET_DATA  => dm9000a_ENET_DATA,                                                          --                      .export
			ENET_CMD   => dm9000a_ENET_CMD,                                                           --                      .export
			ENET_RD_N  => dm9000a_ENET_RD_N,                                                          --                      .export
			ENET_WR_N  => dm9000a_ENET_WR_N,                                                          --                      .export
			ENET_CS_N  => dm9000a_ENET_CS_N,                                                          --                      .export
			ENET_RST_N => dm9000a_ENET_RST_N,                                                         --                      .export
			ENET_CLK   => dm9000a_ENET_CLK,                                                           --                      .export
			ENET_INT   => dm9000a_ENET_INT,                                                           --                      .export
			iDATA      => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_writedata,            --        avalon_slave_0.writedata
			iCMD       => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_address(0),           --                      .address
			iRD_N      => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read_ports_inv,       --                      .read_n
			iWR_N      => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write_ports_inv,      --                      .write_n
			iCS_N      => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect_ports_inv, --                      .chipselect_n
			oDATA      => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_readdata,             --                      .readdata
			oINT       => irq_mapper_receiver15_irq                                                   --    avalon_slave_0_irq.irq
		);

	pio_async_reset : component NIOSIImicro_pio_en_mux
		port map (
			clk        => pll_c0_clk,                                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                          --               reset.reset_n
			address    => pio_async_reset_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_async_reset_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_async_reset_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_async_reset_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_async_reset_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pio_async_reset_export                                             -- external_connection.export
		);

	cpu_instruction_master_translator : component niosiimicro_cpu_instruction_master_translator
		generic map (
			AV_ADDRESS_W                => 25,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 25,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 1,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                            --                     reset.reset
			uav_address              => cpu_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read                  => cpu_instruction_master_read,                                               --                          .read
			av_readdata              => cpu_instruction_master_readdata,                                           --                          .readdata
			av_readdatavalid         => cpu_instruction_master_readdatavalid,                                      --                          .readdatavalid
			av_burstcount            => "1",                                                                       --               (terminated)
			av_byteenable            => "1111",                                                                    --               (terminated)
			av_beginbursttransfer    => '0',                                                                       --               (terminated)
			av_begintransfer         => '0',                                                                       --               (terminated)
			av_chipselect            => '0',                                                                       --               (terminated)
			av_write                 => '0',                                                                       --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                        --               (terminated)
			av_lock                  => '0',                                                                       --               (terminated)
			av_debugaccess           => '0',                                                                       --               (terminated)
			uav_clken                => open,                                                                      --               (terminated)
			av_clken                 => '1',                                                                       --               (terminated)
			uav_response             => "00",                                                                      --               (terminated)
			av_response              => open,                                                                      --               (terminated)
			uav_writeresponserequest => open,                                                                      --               (terminated)
			uav_writeresponsevalid   => '0',                                                                       --               (terminated)
			av_writeresponserequest  => '0',                                                                       --               (terminated)
			av_writeresponsevalid    => open                                                                       --               (terminated)
		);

	cpu_data_master_translator : component niosiimicro_cpu_data_master_translator
		generic map (
			AV_ADDRESS_W                => 25,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 25,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 1
		)
		port map (
			clk                      => pll_c0_clk,                                                         --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                     --                     reset.reset
			uav_address              => cpu_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_data_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => cpu_data_master_byteenable,                                         --                          .byteenable
			av_read                  => cpu_data_master_read,                                               --                          .read
			av_readdata              => cpu_data_master_readdata,                                           --                          .readdata
			av_write                 => cpu_data_master_write,                                              --                          .write
			av_writedata             => cpu_data_master_writedata,                                          --                          .writedata
			av_debugaccess           => cpu_data_master_debugaccess,                                        --                          .debugaccess
			av_burstcount            => "1",                                                                --               (terminated)
			av_beginbursttransfer    => '0',                                                                --               (terminated)
			av_begintransfer         => '0',                                                                --               (terminated)
			av_chipselect            => '0',                                                                --               (terminated)
			av_readdatavalid         => open,                                                               --               (terminated)
			av_lock                  => '0',                                                                --               (terminated)
			uav_clken                => open,                                                               --               (terminated)
			av_clken                 => '1',                                                                --               (terminated)
			uav_response             => "00",                                                               --               (terminated)
			av_response              => open,                                                               --               (terminated)
			uav_writeresponserequest => open,                                                               --               (terminated)
			uav_writeresponsevalid   => '0',                                                                --               (terminated)
			av_writeresponserequest  => '0',                                                                --               (terminated)
			av_writeresponsevalid    => open                                                                --               (terminated)
		);

	cpu_jtag_debug_module_translator : component niosiimicro_cpu_jtag_debug_module_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                       --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                   --                    reset.reset
			uav_address              => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => cpu_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => cpu_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => cpu_jtag_debug_module_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                                             --              (terminated)
			av_burstcount            => open,                                                                             --              (terminated)
			av_readdatavalid         => '0',                                                                              --              (terminated)
			av_writebyteenable       => open,                                                                             --              (terminated)
			av_lock                  => open,                                                                             --              (terminated)
			av_chipselect            => open,                                                                             --              (terminated)
			av_clken                 => open,                                                                             --              (terminated)
			uav_clken                => '0',                                                                              --              (terminated)
			av_outputenable          => open,                                                                             --              (terminated)
			uav_response             => open,                                                                             --              (terminated)
			av_response              => "00",                                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                                             --              (terminated)
			av_writeresponserequest  => open,                                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                                               --              (terminated)
		);

	sdram_s1_translator : component niosiimicro_sdram_s1_translator
		generic map (
			AV_ADDRESS_W                   => 22,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                          --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                      --                    reset.reset
			uav_address              => sdram_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sdram_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sdram_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sdram_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sdram_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => sdram_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => sdram_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sdram_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => sdram_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => sdram_s1_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => sdram_s1_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => sdram_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                --              (terminated)
			av_beginbursttransfer    => open,                                                                --              (terminated)
			av_burstcount            => open,                                                                --              (terminated)
			av_writebyteenable       => open,                                                                --              (terminated)
			av_lock                  => open,                                                                --              (terminated)
			av_clken                 => open,                                                                --              (terminated)
			uav_clken                => '0',                                                                 --              (terminated)
			av_debugaccess           => open,                                                                --              (terminated)
			av_outputenable          => open,                                                                --              (terminated)
			uav_response             => open,                                                                --              (terminated)
			av_response              => "00",                                                                --              (terminated)
			uav_writeresponserequest => '0',                                                                 --              (terminated)
			uav_writeresponsevalid   => open,                                                                --              (terminated)
			av_writeresponserequest  => open,                                                                --              (terminated)
			av_writeresponsevalid    => '0'                                                                  --              (terminated)
		);

	system_id_control_slave_translator : component niosiimicro_system_id_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                         --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                     --                    reset.reset
			uav_address              => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => system_id_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => system_id_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                               --              (terminated)
			av_read                  => open,                                                                               --              (terminated)
			av_writedata             => open,                                                                               --              (terminated)
			av_begintransfer         => open,                                                                               --              (terminated)
			av_beginbursttransfer    => open,                                                                               --              (terminated)
			av_burstcount            => open,                                                                               --              (terminated)
			av_byteenable            => open,                                                                               --              (terminated)
			av_readdatavalid         => '0',                                                                                --              (terminated)
			av_waitrequest           => '0',                                                                                --              (terminated)
			av_writebyteenable       => open,                                                                               --              (terminated)
			av_lock                  => open,                                                                               --              (terminated)
			av_chipselect            => open,                                                                               --              (terminated)
			av_clken                 => open,                                                                               --              (terminated)
			uav_clken                => '0',                                                                                --              (terminated)
			av_debugaccess           => open,                                                                               --              (terminated)
			av_outputenable          => open,                                                                               --              (terminated)
			uav_response             => open,                                                                               --              (terminated)
			av_response              => "00",                                                                               --              (terminated)
			uav_writeresponserequest => '0',                                                                                --              (terminated)
			uav_writeresponsevalid   => open,                                                                               --              (terminated)
			av_writeresponserequest  => open,                                                                               --              (terminated)
			av_writeresponsevalid    => '0'                                                                                 --              (terminated)
		);

	pll_pll_slave_translator : component niosiimicro_pll_pll_slave_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50_clk,                                                               --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                       --                    reset.reset
			uav_address              => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pll_pll_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pll_pll_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => pll_pll_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => pll_pll_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pll_pll_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer         => open,                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                     --              (terminated)
			av_burstcount            => open,                                                                     --              (terminated)
			av_byteenable            => open,                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                      --              (terminated)
			av_waitrequest           => '0',                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                     --              (terminated)
			av_lock                  => open,                                                                     --              (terminated)
			av_chipselect            => open,                                                                     --              (terminated)
			av_clken                 => open,                                                                     --              (terminated)
			uav_clken                => '0',                                                                      --              (terminated)
			av_debugaccess           => open,                                                                     --              (terminated)
			av_outputenable          => open,                                                                     --              (terminated)
			uav_response             => open,                                                                     --              (terminated)
			av_response              => "00",                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                       --              (terminated)
		);

	uart_avalon_jtag_slave_translator : component niosiimicro_uart_avalon_jtag_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                        --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                    --                    reset.reset
			uav_address              => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                                              --              (terminated)
			av_burstcount            => open,                                                                              --              (terminated)
			av_byteenable            => open,                                                                              --              (terminated)
			av_readdatavalid         => '0',                                                                               --              (terminated)
			av_writebyteenable       => open,                                                                              --              (terminated)
			av_lock                  => open,                                                                              --              (terminated)
			av_clken                 => open,                                                                              --              (terminated)
			uav_clken                => '0',                                                                               --              (terminated)
			av_debugaccess           => open,                                                                              --              (terminated)
			av_outputenable          => open,                                                                              --              (terminated)
			uav_response             => open,                                                                              --              (terminated)
			av_response              => "00",                                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                                              --              (terminated)
			av_writeresponserequest  => open,                                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                                --              (terminated)
		);

	timer_0_s1_translator : component niosiimicro_timer_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                            --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => timer_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => timer_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => timer_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => timer_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => timer_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	timer_1_s1_translator : component niosiimicro_timer_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                            --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => timer_1_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => timer_1_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => timer_1_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => timer_1_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => timer_1_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	pio_in_sw_s1_translator : component niosiimicro_pio_in_sw_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                              --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                          --                    reset.reset
			uav_address              => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_in_sw_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => pio_in_sw_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                    --              (terminated)
			av_read                  => open,                                                                    --              (terminated)
			av_writedata             => open,                                                                    --              (terminated)
			av_begintransfer         => open,                                                                    --              (terminated)
			av_beginbursttransfer    => open,                                                                    --              (terminated)
			av_burstcount            => open,                                                                    --              (terminated)
			av_byteenable            => open,                                                                    --              (terminated)
			av_readdatavalid         => '0',                                                                     --              (terminated)
			av_waitrequest           => '0',                                                                     --              (terminated)
			av_writebyteenable       => open,                                                                    --              (terminated)
			av_lock                  => open,                                                                    --              (terminated)
			av_chipselect            => open,                                                                    --              (terminated)
			av_clken                 => open,                                                                    --              (terminated)
			uav_clken                => '0',                                                                     --              (terminated)
			av_debugaccess           => open,                                                                    --              (terminated)
			av_outputenable          => open,                                                                    --              (terminated)
			uav_response             => open,                                                                    --              (terminated)
			av_response              => "00",                                                                    --              (terminated)
			uav_writeresponserequest => '0',                                                                     --              (terminated)
			uav_writeresponsevalid   => open,                                                                    --              (terminated)
			av_writeresponserequest  => open,                                                                    --              (terminated)
			av_writeresponsevalid    => '0'                                                                      --              (terminated)
		);

	pio_in_key_edge_s1_translator : component niosiimicro_pio_in_key_edge_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                    --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                --                    reset.reset
			uav_address              => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_in_key_edge_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_in_key_edge_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_in_key_edge_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_in_key_edge_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_in_key_edge_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                          --              (terminated)
			av_begintransfer         => open,                                                                          --              (terminated)
			av_beginbursttransfer    => open,                                                                          --              (terminated)
			av_burstcount            => open,                                                                          --              (terminated)
			av_byteenable            => open,                                                                          --              (terminated)
			av_readdatavalid         => '0',                                                                           --              (terminated)
			av_waitrequest           => '0',                                                                           --              (terminated)
			av_writebyteenable       => open,                                                                          --              (terminated)
			av_lock                  => open,                                                                          --              (terminated)
			av_clken                 => open,                                                                          --              (terminated)
			uav_clken                => '0',                                                                           --              (terminated)
			av_debugaccess           => open,                                                                          --              (terminated)
			av_outputenable          => open,                                                                          --              (terminated)
			uav_response             => open,                                                                          --              (terminated)
			av_response              => "00",                                                                          --              (terminated)
			uav_writeresponserequest => '0',                                                                           --              (terminated)
			uav_writeresponsevalid   => open,                                                                          --              (terminated)
			av_writeresponserequest  => open,                                                                          --              (terminated)
			av_writeresponsevalid    => '0'                                                                            --              (terminated)
		);

	pio_in_ext_s1_translator : component niosiimicro_pio_in_key_edge_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                           --                    reset.reset
			uav_address              => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_in_ext_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_in_ext_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_in_ext_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_in_ext_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_in_ext_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                     --              (terminated)
			av_begintransfer         => open,                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                     --              (terminated)
			av_burstcount            => open,                                                                     --              (terminated)
			av_byteenable            => open,                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                      --              (terminated)
			av_waitrequest           => '0',                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                     --              (terminated)
			av_lock                  => open,                                                                     --              (terminated)
			av_clken                 => open,                                                                     --              (terminated)
			uav_clken                => '0',                                                                      --              (terminated)
			av_debugaccess           => open,                                                                     --              (terminated)
			av_outputenable          => open,                                                                     --              (terminated)
			uav_response             => open,                                                                     --              (terminated)
			av_response              => "00",                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                       --              (terminated)
		);

	pio_out_red_s1_translator : component niosiimicro_pio_out_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                            --                    reset.reset
			uav_address              => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_out_red_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_out_red_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_out_red_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_out_red_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_out_red_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                      --              (terminated)
			av_begintransfer         => open,                                                                      --              (terminated)
			av_beginbursttransfer    => open,                                                                      --              (terminated)
			av_burstcount            => open,                                                                      --              (terminated)
			av_byteenable            => open,                                                                      --              (terminated)
			av_readdatavalid         => '0',                                                                       --              (terminated)
			av_waitrequest           => '0',                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                      --              (terminated)
			av_lock                  => open,                                                                      --              (terminated)
			av_clken                 => open,                                                                      --              (terminated)
			uav_clken                => '0',                                                                       --              (terminated)
			av_debugaccess           => open,                                                                      --              (terminated)
			av_outputenable          => open,                                                                      --              (terminated)
			uav_response             => open,                                                                      --              (terminated)
			av_response              => "00",                                                                      --              (terminated)
			uav_writeresponserequest => '0',                                                                       --              (terminated)
			uav_writeresponsevalid   => open,                                                                      --              (terminated)
			av_writeresponserequest  => open,                                                                      --              (terminated)
			av_writeresponsevalid    => '0'                                                                        --              (terminated)
		);

	pio_out_green_s1_translator : component niosiimicro_pio_out_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                  --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                              --                    reset.reset
			uav_address              => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_out_green_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_out_green_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_out_green_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_out_green_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_out_green_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                        --              (terminated)
			av_begintransfer         => open,                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                        --              (terminated)
			av_burstcount            => open,                                                                        --              (terminated)
			av_byteenable            => open,                                                                        --              (terminated)
			av_readdatavalid         => '0',                                                                         --              (terminated)
			av_waitrequest           => '0',                                                                         --              (terminated)
			av_writebyteenable       => open,                                                                        --              (terminated)
			av_lock                  => open,                                                                        --              (terminated)
			av_clken                 => open,                                                                        --              (terminated)
			uav_clken                => '0',                                                                         --              (terminated)
			av_debugaccess           => open,                                                                        --              (terminated)
			av_outputenable          => open,                                                                        --              (terminated)
			uav_response             => open,                                                                        --              (terminated)
			av_response              => "00",                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                          --              (terminated)
		);

	pio_out_ext_s1_translator : component niosiimicro_pio_out_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                            --                    reset.reset
			uav_address              => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_out_ext_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_out_ext_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_out_ext_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_out_ext_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_out_ext_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                      --              (terminated)
			av_begintransfer         => open,                                                                      --              (terminated)
			av_beginbursttransfer    => open,                                                                      --              (terminated)
			av_burstcount            => open,                                                                      --              (terminated)
			av_byteenable            => open,                                                                      --              (terminated)
			av_readdatavalid         => '0',                                                                       --              (terminated)
			av_waitrequest           => '0',                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                      --              (terminated)
			av_lock                  => open,                                                                      --              (terminated)
			av_clken                 => open,                                                                      --              (terminated)
			uav_clken                => '0',                                                                       --              (terminated)
			av_debugaccess           => open,                                                                      --              (terminated)
			av_outputenable          => open,                                                                      --              (terminated)
			uav_response             => open,                                                                      --              (terminated)
			av_response              => "00",                                                                      --              (terminated)
			uav_writeresponserequest => '0',                                                                       --              (terminated)
			uav_writeresponsevalid   => open,                                                                      --              (terminated)
			av_writeresponserequest  => open,                                                                      --              (terminated)
			av_writeresponsevalid    => '0'                                                                        --              (terminated)
		);

	pio_async_reset_s1_translator : component niosiimicro_pio_out_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                    --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                --                    reset.reset
			uav_address              => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_async_reset_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_async_reset_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_async_reset_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_async_reset_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_async_reset_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                          --              (terminated)
			av_begintransfer         => open,                                                                          --              (terminated)
			av_beginbursttransfer    => open,                                                                          --              (terminated)
			av_burstcount            => open,                                                                          --              (terminated)
			av_byteenable            => open,                                                                          --              (terminated)
			av_readdatavalid         => '0',                                                                           --              (terminated)
			av_waitrequest           => '0',                                                                           --              (terminated)
			av_writebyteenable       => open,                                                                          --              (terminated)
			av_lock                  => open,                                                                          --              (terminated)
			av_clken                 => open,                                                                          --              (terminated)
			uav_clken                => '0',                                                                           --              (terminated)
			av_debugaccess           => open,                                                                          --              (terminated)
			av_outputenable          => open,                                                                          --              (terminated)
			uav_response             => open,                                                                          --              (terminated)
			av_response              => "00",                                                                          --              (terminated)
			uav_writeresponserequest => '0',                                                                           --              (terminated)
			uav_writeresponsevalid   => open,                                                                          --              (terminated)
			av_writeresponserequest  => open,                                                                          --              (terminated)
			av_writeresponsevalid    => '0'                                                                            --              (terminated)
		);

	pio_en_mux_s1_translator : component niosiimicro_pio_out_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                           --                    reset.reset
			uav_address              => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_en_mux_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_en_mux_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_en_mux_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_en_mux_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_en_mux_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                     --              (terminated)
			av_begintransfer         => open,                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                     --              (terminated)
			av_burstcount            => open,                                                                     --              (terminated)
			av_byteenable            => open,                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                      --              (terminated)
			av_waitrequest           => '0',                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                     --              (terminated)
			av_lock                  => open,                                                                     --              (terminated)
			av_clken                 => open,                                                                     --              (terminated)
			uav_clken                => '0',                                                                      --              (terminated)
			av_debugaccess           => open,                                                                     --              (terminated)
			av_outputenable          => open,                                                                     --              (terminated)
			uav_response             => open,                                                                     --              (terminated)
			av_response              => "00",                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                       --              (terminated)
		);

	pio_direc_s1_translator : component niosiimicro_pio_out_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                              --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                          --                    reset.reset
			uav_address              => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_direc_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_direc_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_direc_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_direc_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_direc_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                    --              (terminated)
			av_begintransfer         => open,                                                                    --              (terminated)
			av_beginbursttransfer    => open,                                                                    --              (terminated)
			av_burstcount            => open,                                                                    --              (terminated)
			av_byteenable            => open,                                                                    --              (terminated)
			av_readdatavalid         => '0',                                                                     --              (terminated)
			av_waitrequest           => '0',                                                                     --              (terminated)
			av_writebyteenable       => open,                                                                    --              (terminated)
			av_lock                  => open,                                                                    --              (terminated)
			av_clken                 => open,                                                                    --              (terminated)
			uav_clken                => '0',                                                                     --              (terminated)
			av_debugaccess           => open,                                                                    --              (terminated)
			av_outputenable          => open,                                                                    --              (terminated)
			uav_response             => open,                                                                    --              (terminated)
			av_response              => "00",                                                                    --              (terminated)
			uav_writeresponserequest => '0',                                                                     --              (terminated)
			uav_writeresponsevalid   => open,                                                                    --              (terminated)
			av_writeresponserequest  => open,                                                                    --              (terminated)
			av_writeresponsevalid    => '0'                                                                      --              (terminated)
		);

	pio_direc_ram_s1_translator : component niosiimicro_pio_out_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                  --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                              --                    reset.reset
			uav_address              => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_direc_ram_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_direc_ram_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_direc_ram_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_direc_ram_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_direc_ram_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                        --              (terminated)
			av_begintransfer         => open,                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                        --              (terminated)
			av_burstcount            => open,                                                                        --              (terminated)
			av_byteenable            => open,                                                                        --              (terminated)
			av_readdatavalid         => '0',                                                                         --              (terminated)
			av_waitrequest           => '0',                                                                         --              (terminated)
			av_writebyteenable       => open,                                                                        --              (terminated)
			av_lock                  => open,                                                                        --              (terminated)
			av_clken                 => open,                                                                        --              (terminated)
			uav_clken                => '0',                                                                         --              (terminated)
			av_debugaccess           => open,                                                                        --              (terminated)
			av_outputenable          => open,                                                                        --              (terminated)
			uav_response             => open,                                                                        --              (terminated)
			av_response              => "00",                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                          --              (terminated)
		);

	pio_wr_s1_translator : component niosiimicro_pio_out_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                           --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                       --                    reset.reset
			uav_address              => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_wr_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_wr_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_wr_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_wr_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_wr_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                 --              (terminated)
			av_begintransfer         => open,                                                                 --              (terminated)
			av_beginbursttransfer    => open,                                                                 --              (terminated)
			av_burstcount            => open,                                                                 --              (terminated)
			av_byteenable            => open,                                                                 --              (terminated)
			av_readdatavalid         => '0',                                                                  --              (terminated)
			av_waitrequest           => '0',                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                 --              (terminated)
			av_lock                  => open,                                                                 --              (terminated)
			av_clken                 => open,                                                                 --              (terminated)
			uav_clken                => '0',                                                                  --              (terminated)
			av_debugaccess           => open,                                                                 --              (terminated)
			av_outputenable          => open,                                                                 --              (terminated)
			uav_response             => open,                                                                 --              (terminated)
			av_response              => "00",                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                   --              (terminated)
		);

	pio_sel_salida_s1_translator : component niosiimicro_pio_out_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                   --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                               --                    reset.reset
			uav_address              => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_sel_salida_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_sel_salida_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_sel_salida_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_sel_salida_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_sel_salida_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                         --              (terminated)
			av_begintransfer         => open,                                                                         --              (terminated)
			av_beginbursttransfer    => open,                                                                         --              (terminated)
			av_burstcount            => open,                                                                         --              (terminated)
			av_byteenable            => open,                                                                         --              (terminated)
			av_readdatavalid         => '0',                                                                          --              (terminated)
			av_waitrequest           => '0',                                                                          --              (terminated)
			av_writebyteenable       => open,                                                                         --              (terminated)
			av_lock                  => open,                                                                         --              (terminated)
			av_clken                 => open,                                                                         --              (terminated)
			uav_clken                => '0',                                                                          --              (terminated)
			av_debugaccess           => open,                                                                         --              (terminated)
			av_outputenable          => open,                                                                         --              (terminated)
			uav_response             => open,                                                                         --              (terminated)
			av_response              => "00",                                                                         --              (terminated)
			uav_writeresponserequest => '0',                                                                          --              (terminated)
			uav_writeresponsevalid   => open,                                                                         --              (terminated)
			av_writeresponserequest  => open,                                                                         --              (terminated)
			av_writeresponsevalid    => '0'                                                                           --              (terminated)
		);

	pio_datos_s1_translator : component niosiimicro_pio_out_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                              --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                          --                    reset.reset
			uav_address              => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_datos_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_datos_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_datos_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_datos_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_datos_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                    --              (terminated)
			av_begintransfer         => open,                                                                    --              (terminated)
			av_beginbursttransfer    => open,                                                                    --              (terminated)
			av_burstcount            => open,                                                                    --              (terminated)
			av_byteenable            => open,                                                                    --              (terminated)
			av_readdatavalid         => '0',                                                                     --              (terminated)
			av_waitrequest           => '0',                                                                     --              (terminated)
			av_writebyteenable       => open,                                                                    --              (terminated)
			av_lock                  => open,                                                                    --              (terminated)
			av_clken                 => open,                                                                    --              (terminated)
			uav_clken                => '0',                                                                     --              (terminated)
			av_debugaccess           => open,                                                                    --              (terminated)
			av_outputenable          => open,                                                                    --              (terminated)
			uav_response             => open,                                                                    --              (terminated)
			av_response              => "00",                                                                    --              (terminated)
			uav_writeresponserequest => '0',                                                                     --              (terminated)
			uav_writeresponsevalid   => open,                                                                    --              (terminated)
			av_writeresponserequest  => open,                                                                    --              (terminated)
			av_writeresponsevalid    => '0'                                                                      --              (terminated)
		);

	pio_compara_int_0_s1_translator : component niosiimicro_pio_in_key_edge_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                      --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                  --                    reset.reset
			uav_address              => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_compara_int_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_compara_int_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_compara_int_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_compara_int_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_compara_int_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                            --              (terminated)
			av_begintransfer         => open,                                                                            --              (terminated)
			av_beginbursttransfer    => open,                                                                            --              (terminated)
			av_burstcount            => open,                                                                            --              (terminated)
			av_byteenable            => open,                                                                            --              (terminated)
			av_readdatavalid         => '0',                                                                             --              (terminated)
			av_waitrequest           => '0',                                                                             --              (terminated)
			av_writebyteenable       => open,                                                                            --              (terminated)
			av_lock                  => open,                                                                            --              (terminated)
			av_clken                 => open,                                                                            --              (terminated)
			uav_clken                => '0',                                                                             --              (terminated)
			av_debugaccess           => open,                                                                            --              (terminated)
			av_outputenable          => open,                                                                            --              (terminated)
			uav_response             => open,                                                                            --              (terminated)
			av_response              => "00",                                                                            --              (terminated)
			uav_writeresponserequest => '0',                                                                             --              (terminated)
			uav_writeresponsevalid   => open,                                                                            --              (terminated)
			av_writeresponserequest  => open,                                                                            --              (terminated)
			av_writeresponsevalid    => '0'                                                                              --              (terminated)
		);

	pio_compara_int_1_s1_translator : component niosiimicro_pio_in_key_edge_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                      --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                  --                    reset.reset
			uav_address              => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_compara_int_1_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_compara_int_1_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_compara_int_1_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_compara_int_1_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_compara_int_1_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                            --              (terminated)
			av_begintransfer         => open,                                                                            --              (terminated)
			av_beginbursttransfer    => open,                                                                            --              (terminated)
			av_burstcount            => open,                                                                            --              (terminated)
			av_byteenable            => open,                                                                            --              (terminated)
			av_readdatavalid         => '0',                                                                             --              (terminated)
			av_waitrequest           => '0',                                                                             --              (terminated)
			av_writebyteenable       => open,                                                                            --              (terminated)
			av_lock                  => open,                                                                            --              (terminated)
			av_clken                 => open,                                                                            --              (terminated)
			uav_clken                => '0',                                                                             --              (terminated)
			av_debugaccess           => open,                                                                            --              (terminated)
			av_outputenable          => open,                                                                            --              (terminated)
			uav_response             => open,                                                                            --              (terminated)
			av_response              => "00",                                                                            --              (terminated)
			uav_writeresponserequest => '0',                                                                             --              (terminated)
			uav_writeresponsevalid   => open,                                                                            --              (terminated)
			av_writeresponserequest  => open,                                                                            --              (terminated)
			av_writeresponsevalid    => '0'                                                                              --              (terminated)
		);

	pio_compara_int_2_s1_translator : component niosiimicro_pio_in_key_edge_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                      --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                  --                    reset.reset
			uav_address              => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_compara_int_2_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_compara_int_2_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_compara_int_2_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_compara_int_2_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_compara_int_2_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                            --              (terminated)
			av_begintransfer         => open,                                                                            --              (terminated)
			av_beginbursttransfer    => open,                                                                            --              (terminated)
			av_burstcount            => open,                                                                            --              (terminated)
			av_byteenable            => open,                                                                            --              (terminated)
			av_readdatavalid         => '0',                                                                             --              (terminated)
			av_waitrequest           => '0',                                                                             --              (terminated)
			av_writebyteenable       => open,                                                                            --              (terminated)
			av_lock                  => open,                                                                            --              (terminated)
			av_clken                 => open,                                                                            --              (terminated)
			uav_clken                => '0',                                                                             --              (terminated)
			av_debugaccess           => open,                                                                            --              (terminated)
			av_outputenable          => open,                                                                            --              (terminated)
			uav_response             => open,                                                                            --              (terminated)
			av_response              => "00",                                                                            --              (terminated)
			uav_writeresponserequest => '0',                                                                             --              (terminated)
			uav_writeresponsevalid   => open,                                                                            --              (terminated)
			av_writeresponserequest  => open,                                                                            --              (terminated)
			av_writeresponsevalid    => '0'                                                                              --              (terminated)
		);

	pio_compara_int_3_s1_translator : component niosiimicro_pio_in_key_edge_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                      --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                  --                    reset.reset
			uav_address              => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_compara_int_3_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_compara_int_3_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_compara_int_3_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_compara_int_3_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_compara_int_3_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                            --              (terminated)
			av_begintransfer         => open,                                                                            --              (terminated)
			av_beginbursttransfer    => open,                                                                            --              (terminated)
			av_burstcount            => open,                                                                            --              (terminated)
			av_byteenable            => open,                                                                            --              (terminated)
			av_readdatavalid         => '0',                                                                             --              (terminated)
			av_waitrequest           => '0',                                                                             --              (terminated)
			av_writebyteenable       => open,                                                                            --              (terminated)
			av_lock                  => open,                                                                            --              (terminated)
			av_clken                 => open,                                                                            --              (terminated)
			uav_clken                => '0',                                                                             --              (terminated)
			av_debugaccess           => open,                                                                            --              (terminated)
			av_outputenable          => open,                                                                            --              (terminated)
			uav_response             => open,                                                                            --              (terminated)
			av_response              => "00",                                                                            --              (terminated)
			uav_writeresponserequest => '0',                                                                             --              (terminated)
			uav_writeresponsevalid   => open,                                                                            --              (terminated)
			av_writeresponserequest  => open,                                                                            --              (terminated)
			av_writeresponsevalid    => '0'                                                                              --              (terminated)
		);

	pio_compara_int_4_s1_translator : component niosiimicro_pio_in_key_edge_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                      --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                  --                    reset.reset
			uav_address              => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_compara_int_4_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_compara_int_4_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_compara_int_4_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_compara_int_4_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_compara_int_4_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                            --              (terminated)
			av_begintransfer         => open,                                                                            --              (terminated)
			av_beginbursttransfer    => open,                                                                            --              (terminated)
			av_burstcount            => open,                                                                            --              (terminated)
			av_byteenable            => open,                                                                            --              (terminated)
			av_readdatavalid         => '0',                                                                             --              (terminated)
			av_waitrequest           => '0',                                                                             --              (terminated)
			av_writebyteenable       => open,                                                                            --              (terminated)
			av_lock                  => open,                                                                            --              (terminated)
			av_clken                 => open,                                                                            --              (terminated)
			uav_clken                => '0',                                                                             --              (terminated)
			av_debugaccess           => open,                                                                            --              (terminated)
			av_outputenable          => open,                                                                            --              (terminated)
			uav_response             => open,                                                                            --              (terminated)
			av_response              => "00",                                                                            --              (terminated)
			uav_writeresponserequest => '0',                                                                             --              (terminated)
			uav_writeresponsevalid   => open,                                                                            --              (terminated)
			av_writeresponserequest  => open,                                                                            --              (terminated)
			av_writeresponsevalid    => '0'                                                                              --              (terminated)
		);

	pio_captura_0_s1_translator : component niosiimicro_pio_in_key_edge_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                  --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                              --                    reset.reset
			uav_address              => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_captura_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_captura_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_captura_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_captura_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_captura_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                        --              (terminated)
			av_begintransfer         => open,                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                        --              (terminated)
			av_burstcount            => open,                                                                        --              (terminated)
			av_byteenable            => open,                                                                        --              (terminated)
			av_readdatavalid         => '0',                                                                         --              (terminated)
			av_waitrequest           => '0',                                                                         --              (terminated)
			av_writebyteenable       => open,                                                                        --              (terminated)
			av_lock                  => open,                                                                        --              (terminated)
			av_clken                 => open,                                                                        --              (terminated)
			uav_clken                => '0',                                                                         --              (terminated)
			av_debugaccess           => open,                                                                        --              (terminated)
			av_outputenable          => open,                                                                        --              (terminated)
			uav_response             => open,                                                                        --              (terminated)
			av_response              => "00",                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                          --              (terminated)
		);

	pio_captura_1_s1_translator : component niosiimicro_pio_in_key_edge_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                  --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                              --                    reset.reset
			uav_address              => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_captura_1_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_captura_1_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_captura_1_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_captura_1_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_captura_1_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                        --              (terminated)
			av_begintransfer         => open,                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                        --              (terminated)
			av_burstcount            => open,                                                                        --              (terminated)
			av_byteenable            => open,                                                                        --              (terminated)
			av_readdatavalid         => '0',                                                                         --              (terminated)
			av_waitrequest           => '0',                                                                         --              (terminated)
			av_writebyteenable       => open,                                                                        --              (terminated)
			av_lock                  => open,                                                                        --              (terminated)
			av_clken                 => open,                                                                        --              (terminated)
			uav_clken                => '0',                                                                         --              (terminated)
			av_debugaccess           => open,                                                                        --              (terminated)
			av_outputenable          => open,                                                                        --              (terminated)
			uav_response             => open,                                                                        --              (terminated)
			av_response              => "00",                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                          --              (terminated)
		);

	pio_captura_2_s1_translator : component niosiimicro_pio_in_key_edge_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                  --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                              --                    reset.reset
			uav_address              => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_captura_2_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_captura_2_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_captura_2_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_captura_2_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_captura_2_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                        --              (terminated)
			av_begintransfer         => open,                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                        --              (terminated)
			av_burstcount            => open,                                                                        --              (terminated)
			av_byteenable            => open,                                                                        --              (terminated)
			av_readdatavalid         => '0',                                                                         --              (terminated)
			av_waitrequest           => '0',                                                                         --              (terminated)
			av_writebyteenable       => open,                                                                        --              (terminated)
			av_lock                  => open,                                                                        --              (terminated)
			av_clken                 => open,                                                                        --              (terminated)
			uav_clken                => '0',                                                                         --              (terminated)
			av_debugaccess           => open,                                                                        --              (terminated)
			av_outputenable          => open,                                                                        --              (terminated)
			uav_response             => open,                                                                        --              (terminated)
			av_response              => "00",                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                          --              (terminated)
		);

	pio_captura_3_s1_translator : component niosiimicro_pio_in_key_edge_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                  --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                              --                    reset.reset
			uav_address              => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_captura_3_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_captura_3_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_captura_3_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_captura_3_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_captura_3_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                        --              (terminated)
			av_begintransfer         => open,                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                        --              (terminated)
			av_burstcount            => open,                                                                        --              (terminated)
			av_byteenable            => open,                                                                        --              (terminated)
			av_readdatavalid         => '0',                                                                         --              (terminated)
			av_waitrequest           => '0',                                                                         --              (terminated)
			av_writebyteenable       => open,                                                                        --              (terminated)
			av_lock                  => open,                                                                        --              (terminated)
			av_clken                 => open,                                                                        --              (terminated)
			uav_clken                => '0',                                                                         --              (terminated)
			av_debugaccess           => open,                                                                        --              (terminated)
			av_outputenable          => open,                                                                        --              (terminated)
			uav_response             => open,                                                                        --              (terminated)
			av_response              => "00",                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                          --              (terminated)
		);

	pio_captura_4_s1_translator : component niosiimicro_pio_in_key_edge_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                  --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                              --                    reset.reset
			uav_address              => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_captura_4_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_captura_4_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_captura_4_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_captura_4_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_captura_4_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                        --              (terminated)
			av_begintransfer         => open,                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                        --              (terminated)
			av_burstcount            => open,                                                                        --              (terminated)
			av_byteenable            => open,                                                                        --              (terminated)
			av_readdatavalid         => '0',                                                                         --              (terminated)
			av_waitrequest           => '0',                                                                         --              (terminated)
			av_writebyteenable       => open,                                                                        --              (terminated)
			av_lock                  => open,                                                                        --              (terminated)
			av_clken                 => open,                                                                        --              (terminated)
			uav_clken                => '0',                                                                         --              (terminated)
			av_debugaccess           => open,                                                                        --              (terminated)
			av_outputenable          => open,                                                                        --              (terminated)
			uav_response             => open,                                                                        --              (terminated)
			av_response              => "00",                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                          --              (terminated)
		);

	pio_in_32_s1_translator : component niosiimicro_pio_in_key_edge_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                              --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                          --                    reset.reset
			uav_address              => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_in_32_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_in_32_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_in_32_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_in_32_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_in_32_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                    --              (terminated)
			av_begintransfer         => open,                                                                    --              (terminated)
			av_beginbursttransfer    => open,                                                                    --              (terminated)
			av_burstcount            => open,                                                                    --              (terminated)
			av_byteenable            => open,                                                                    --              (terminated)
			av_readdatavalid         => '0',                                                                     --              (terminated)
			av_waitrequest           => '0',                                                                     --              (terminated)
			av_writebyteenable       => open,                                                                    --              (terminated)
			av_lock                  => open,                                                                    --              (terminated)
			av_clken                 => open,                                                                    --              (terminated)
			uav_clken                => '0',                                                                     --              (terminated)
			av_debugaccess           => open,                                                                    --              (terminated)
			av_outputenable          => open,                                                                    --              (terminated)
			uav_response             => open,                                                                    --              (terminated)
			av_response              => "00",                                                                    --              (terminated)
			uav_writeresponserequest => '0',                                                                     --              (terminated)
			uav_writeresponsevalid   => open,                                                                    --              (terminated)
			av_writeresponserequest  => open,                                                                    --              (terminated)
			av_writeresponsevalid    => '0'                                                                      --              (terminated)
		);

	lcd_control_slave_translator : component niosiimicro_lcd_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 8,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 13,
			AV_WRITE_WAIT_CYCLES           => 13,
			AV_SETUP_WAIT_CYCLES           => 13,
			AV_DATA_HOLD_CYCLES            => 13
		)
		port map (
			clk                      => pll_c0_clk,                                                                   --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                               --                    reset.reset
			uav_address              => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => lcd_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => lcd_control_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => lcd_control_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => lcd_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => lcd_control_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer         => lcd_control_slave_translator_avalon_anti_slave_0_begintransfer,               --                         .begintransfer
			av_beginbursttransfer    => open,                                                                         --              (terminated)
			av_burstcount            => open,                                                                         --              (terminated)
			av_byteenable            => open,                                                                         --              (terminated)
			av_readdatavalid         => '0',                                                                          --              (terminated)
			av_waitrequest           => '0',                                                                          --              (terminated)
			av_writebyteenable       => open,                                                                         --              (terminated)
			av_lock                  => open,                                                                         --              (terminated)
			av_chipselect            => open,                                                                         --              (terminated)
			av_clken                 => open,                                                                         --              (terminated)
			uav_clken                => '0',                                                                          --              (terminated)
			av_debugaccess           => open,                                                                         --              (terminated)
			av_outputenable          => open,                                                                         --              (terminated)
			uav_response             => open,                                                                         --              (terminated)
			av_response              => "00",                                                                         --              (terminated)
			uav_writeresponserequest => '0',                                                                          --              (terminated)
			uav_writeresponsevalid   => open,                                                                         --              (terminated)
			av_writeresponserequest  => open,                                                                         --              (terminated)
			av_writeresponsevalid    => '0'                                                                           --              (terminated)
		);

	dm9000a_avalon_slave_0_translator : component niosiimicro_dm9000a_avalon_slave_0_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 2,
			AV_WRITE_WAIT_CYCLES           => 2,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => pll_c0_clk,                                                                        --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                    --                    reset.reset
			uav_address              => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                                              --              (terminated)
			av_burstcount            => open,                                                                              --              (terminated)
			av_byteenable            => open,                                                                              --              (terminated)
			av_readdatavalid         => '0',                                                                               --              (terminated)
			av_waitrequest           => '0',                                                                               --              (terminated)
			av_writebyteenable       => open,                                                                              --              (terminated)
			av_lock                  => open,                                                                              --              (terminated)
			av_clken                 => open,                                                                              --              (terminated)
			uav_clken                => '0',                                                                               --              (terminated)
			av_debugaccess           => open,                                                                              --              (terminated)
			av_outputenable          => open,                                                                              --              (terminated)
			uav_response             => open,                                                                              --              (terminated)
			av_response              => "00",                                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                                              --              (terminated)
			av_writeresponserequest  => open,                                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                                --              (terminated)
		);

	cpu_instruction_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_BEGIN_BURST           => 80,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			PKT_BURST_TYPE_H          => 77,
			PKT_BURST_TYPE_L          => 76,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_TRANS_EXCLUSIVE       => 66,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_THREAD_ID_H           => 94,
			PKT_THREAD_ID_L           => 94,
			PKT_CACHE_H               => 101,
			PKT_CACHE_L               => 98,
			PKT_DATA_SIDEBAND_H       => 79,
			PKT_DATA_SIDEBAND_L       => 79,
			PKT_QOS_H                 => 81,
			PKT_QOS_L                 => 81,
			PKT_ADDR_SIDEBAND_H       => 78,
			PKT_ADDR_SIDEBAND_L       => 78,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			ST_DATA_W                 => 104,
			ST_CHANNEL_W              => 33,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 3,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                         --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			av_address              => cpu_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => limiter_rsp_src_valid,                                                              --        rp.valid
			rp_data                 => limiter_rsp_src_data,                                                               --          .data
			rp_channel              => limiter_rsp_src_channel,                                                            --          .channel
			rp_startofpacket        => limiter_rsp_src_startofpacket,                                                      --          .startofpacket
			rp_endofpacket          => limiter_rsp_src_endofpacket,                                                        --          .endofpacket
			rp_ready                => limiter_rsp_src_ready,                                                              --          .ready
			av_response             => open,                                                                               -- (terminated)
			av_writeresponserequest => '0',                                                                                -- (terminated)
			av_writeresponsevalid   => open                                                                                -- (terminated)
		);

	cpu_data_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_BEGIN_BURST           => 80,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			PKT_BURST_TYPE_H          => 77,
			PKT_BURST_TYPE_L          => 76,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_TRANS_EXCLUSIVE       => 66,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_THREAD_ID_H           => 94,
			PKT_THREAD_ID_L           => 94,
			PKT_CACHE_H               => 101,
			PKT_CACHE_L               => 98,
			PKT_DATA_SIDEBAND_H       => 79,
			PKT_DATA_SIDEBAND_L       => 79,
			PKT_QOS_H                 => 81,
			PKT_QOS_L                 => 81,
			PKT_ADDR_SIDEBAND_H       => 78,
			PKT_ADDR_SIDEBAND_L       => 78,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			ST_DATA_W                 => 104,
			ST_CHANNEL_W              => 33,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                  --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			av_address              => cpu_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_001_src_valid,                                                  --        rp.valid
			rp_data                 => rsp_xbar_mux_001_src_data,                                                   --          .data
			rp_channel              => rsp_xbar_mux_001_src_channel,                                                --          .channel
			rp_startofpacket        => rsp_xbar_mux_001_src_startofpacket,                                          --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_001_src_endofpacket,                                            --          .endofpacket
			rp_ready                => rsp_xbar_mux_001_src_ready,                                                  --          .ready
			av_response             => open,                                                                        -- (terminated)
			av_writeresponserequest => '0',                                                                         -- (terminated)
			av_writeresponsevalid   => open                                                                         -- (terminated)
		);

	cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                                 --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                             --       clk_reset.reset
			m0_address              => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_src_ready,                                                                     --              cp.ready
			cp_valid                => cmd_xbar_mux_src_valid,                                                                     --                .valid
			cp_data                 => cmd_xbar_mux_src_data,                                                                      --                .data
			cp_startofpacket        => cmd_xbar_mux_src_startofpacket,                                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_src_endofpacket,                                                               --                .endofpacket
			cp_channel              => cmd_xbar_mux_src_channel,                                                                   --                .channel
			rf_sink_ready           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                       --     (terminated)
			m0_writeresponserequest => open,                                                                                       --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                         --     (terminated)
		);

	cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                                 --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                             -- clk_reset.reset
			in_data           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                       -- (terminated)
			csr_read          => '0',                                                                                        -- (terminated)
			csr_write         => '0',                                                                                        -- (terminated)
			csr_readdata      => open,                                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                         -- (terminated)
			almost_full_data  => open,                                                                                       -- (terminated)
			almost_empty_data => open,                                                                                       -- (terminated)
			in_empty          => '0',                                                                                        -- (terminated)
			out_empty         => open,                                                                                       -- (terminated)
			in_error          => '0',                                                                                        -- (terminated)
			out_error         => open,                                                                                       -- (terminated)
			in_channel        => '0',                                                                                        -- (terminated)
			out_channel       => open                                                                                        -- (terminated)
		);

	sdram_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_sdram_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 62,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_ADDR_H                => 42,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 43,
			PKT_TRANS_POSTED          => 44,
			PKT_TRANS_WRITE           => 45,
			PKT_TRANS_READ            => 46,
			PKT_TRANS_LOCK            => 47,
			PKT_SRC_ID_H              => 69,
			PKT_SRC_ID_L              => 64,
			PKT_DEST_ID_H             => 75,
			PKT_DEST_ID_L             => 70,
			PKT_BURSTWRAP_H           => 54,
			PKT_BURSTWRAP_L           => 52,
			PKT_BYTE_CNT_H            => 51,
			PKT_BYTE_CNT_L            => 49,
			PKT_PROTECTION_H          => 79,
			PKT_PROTECTION_L          => 77,
			PKT_RESPONSE_STATUS_H     => 85,
			PKT_RESPONSE_STATUS_L     => 84,
			PKT_BURST_SIZE_H          => 57,
			PKT_BURST_SIZE_L          => 55,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 86,
			AVS_BURSTCOUNT_W          => 2,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                    --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                --       clk_reset.reset
			m0_address              => sdram_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sdram_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sdram_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sdram_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_source0_ready,                                                   --              cp.ready
			cp_valid                => burst_adapter_source0_valid,                                                   --                .valid
			cp_data                 => burst_adapter_source0_data,                                                    --                .data
			cp_startofpacket        => burst_adapter_source0_startofpacket,                                           --                .startofpacket
			cp_endofpacket          => burst_adapter_source0_endofpacket,                                             --                .endofpacket
			cp_channel              => burst_adapter_source0_channel,                                                 --                .channel
			rf_sink_ready           => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                          --     (terminated)
			m0_writeresponserequest => open,                                                                          --     (terminated)
			m0_writeresponsevalid   => '0'                                                                            --     (terminated)
		);

	sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 87,
			FIFO_DEPTH          => 8,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                    --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                -- clk_reset.reset
			in_data           => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                          -- (terminated)
			csr_read          => '0',                                                                           -- (terminated)
			csr_write         => '0',                                                                           -- (terminated)
			csr_readdata      => open,                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                            -- (terminated)
			almost_full_data  => open,                                                                          -- (terminated)
			almost_empty_data => open,                                                                          -- (terminated)
			in_empty          => '0',                                                                           -- (terminated)
			out_empty         => open,                                                                          -- (terminated)
			in_error          => '0',                                                                           -- (terminated)
			out_error         => open,                                                                          -- (terminated)
			in_channel        => '0',                                                                           -- (terminated)
			out_channel       => open                                                                           -- (terminated)
		);

	sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component niosiimicro_sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 18,
			FIFO_DEPTH          => 8,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 3,
			USE_MEMORY_BLOCKS   => 1,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                              --       clk.clk
			reset             => rst_controller_reset_out_reset,                                          -- clk_reset.reset
			in_data           => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                    -- (terminated)
			csr_read          => '0',                                                                     -- (terminated)
			csr_write         => '0',                                                                     -- (terminated)
			csr_readdata      => open,                                                                    -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                      -- (terminated)
			almost_full_data  => open,                                                                    -- (terminated)
			almost_empty_data => open,                                                                    -- (terminated)
			in_startofpacket  => '0',                                                                     -- (terminated)
			in_endofpacket    => '0',                                                                     -- (terminated)
			out_startofpacket => open,                                                                    -- (terminated)
			out_endofpacket   => open,                                                                    -- (terminated)
			in_empty          => '0',                                                                     -- (terminated)
			out_empty         => open,                                                                    -- (terminated)
			in_error          => '0',                                                                     -- (terminated)
			out_error         => open,                                                                    -- (terminated)
			in_channel        => '0',                                                                     -- (terminated)
			out_channel       => open                                                                     -- (terminated)
		);

	system_id_control_slave_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                                   --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                               --       clk_reset.reset
			m0_address              => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => system_id_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => system_id_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => system_id_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => system_id_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => system_id_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => system_id_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_002_src_ready,                                                                   --              cp.ready
			cp_valid                => cmd_xbar_mux_002_src_valid,                                                                   --                .valid
			cp_data                 => cmd_xbar_mux_002_src_data,                                                                    --                .data
			cp_startofpacket        => cmd_xbar_mux_002_src_startofpacket,                                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_002_src_endofpacket,                                                             --                .endofpacket
			cp_channel              => cmd_xbar_mux_002_src_channel,                                                                 --                .channel
			rf_sink_ready           => system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => system_id_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => system_id_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => system_id_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => system_id_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => system_id_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => system_id_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => system_id_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => system_id_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => system_id_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => system_id_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => system_id_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                         --     (terminated)
			m0_writeresponserequest => open,                                                                                         --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                           --     (terminated)
		);

	system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                                   --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                               -- clk_reset.reset
			in_data           => system_id_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => system_id_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => system_id_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => system_id_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => system_id_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => system_id_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                         -- (terminated)
			csr_read          => '0',                                                                                          -- (terminated)
			csr_write         => '0',                                                                                          -- (terminated)
			csr_readdata      => open,                                                                                         -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                           -- (terminated)
			almost_full_data  => open,                                                                                         -- (terminated)
			almost_empty_data => open,                                                                                         -- (terminated)
			in_empty          => '0',                                                                                          -- (terminated)
			out_empty         => open,                                                                                         -- (terminated)
			in_error          => '0',                                                                                          -- (terminated)
			out_error         => open,                                                                                         -- (terminated)
			in_channel        => '0',                                                                                          -- (terminated)
			out_channel       => open                                                                                          -- (terminated)
		);

	pll_pll_slave_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50_clk,                                                                         --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                 --       clk_reset.reset
			m0_address              => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => crosser_out_ready,                                                                  --              cp.ready
			cp_valid                => crosser_out_valid,                                                                  --                .valid
			cp_data                 => crosser_out_data,                                                                   --                .data
			cp_startofpacket        => crosser_out_startofpacket,                                                          --                .startofpacket
			cp_endofpacket          => crosser_out_endofpacket,                                                            --                .endofpacket
			cp_channel              => crosser_out_channel,                                                                --                .channel
			rf_sink_ready           => pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                 --     (terminated)
		);

	pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50_clk,                                                                         --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                 -- clk_reset.reset
			in_data           => pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                               -- (terminated)
			csr_read          => '0',                                                                                -- (terminated)
			csr_write         => '0',                                                                                -- (terminated)
			csr_readdata      => open,                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                 -- (terminated)
			almost_full_data  => open,                                                                               -- (terminated)
			almost_empty_data => open,                                                                               -- (terminated)
			in_empty          => '0',                                                                                -- (terminated)
			out_empty         => open,                                                                               -- (terminated)
			in_error          => '0',                                                                                -- (terminated)
			out_error         => open,                                                                               -- (terminated)
			in_channel        => '0',                                                                                -- (terminated)
			out_channel       => open                                                                                -- (terminated)
		);

	pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo : component niosiimicro_pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 34,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50_clk,                                                                   --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                           -- clk_reset.reset
			in_data           => pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                         -- (terminated)
			csr_read          => '0',                                                                          -- (terminated)
			csr_write         => '0',                                                                          -- (terminated)
			csr_readdata      => open,                                                                         -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                           -- (terminated)
			almost_full_data  => open,                                                                         -- (terminated)
			almost_empty_data => open,                                                                         -- (terminated)
			in_startofpacket  => '0',                                                                          -- (terminated)
			in_endofpacket    => '0',                                                                          -- (terminated)
			out_startofpacket => open,                                                                         -- (terminated)
			out_endofpacket   => open,                                                                         -- (terminated)
			in_empty          => '0',                                                                          -- (terminated)
			out_empty         => open,                                                                         -- (terminated)
			in_error          => '0',                                                                          -- (terminated)
			out_error         => open,                                                                         -- (terminated)
			in_channel        => '0',                                                                          -- (terminated)
			out_channel       => open                                                                          -- (terminated)
		);

	uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                                  --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                              --       clk_reset.reset
			m0_address              => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src4_ready,                                                               --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src4_valid,                                                               --                .valid
			cp_data                 => cmd_xbar_demux_001_src4_data,                                                                --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src4_startofpacket,                                                       --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src4_endofpacket,                                                         --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src4_channel,                                                             --                .channel
			rf_sink_ready           => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                          --     (terminated)
		);

	uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                                  --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                              -- clk_reset.reset
			in_data           => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                        -- (terminated)
			csr_read          => '0',                                                                                         -- (terminated)
			csr_write         => '0',                                                                                         -- (terminated)
			csr_readdata      => open,                                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                          -- (terminated)
			almost_full_data  => open,                                                                                        -- (terminated)
			almost_empty_data => open,                                                                                        -- (terminated)
			in_empty          => '0',                                                                                         -- (terminated)
			out_empty         => open,                                                                                        -- (terminated)
			in_error          => '0',                                                                                         -- (terminated)
			out_error         => open,                                                                                        -- (terminated)
			in_channel        => '0',                                                                                         -- (terminated)
			out_channel       => open                                                                                         -- (terminated)
		);

	timer_0_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                      --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src5_ready,                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src5_valid,                                                   --                .valid
			cp_data                 => cmd_xbar_demux_001_src5_data,                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src5_startofpacket,                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src5_endofpacket,                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src5_channel,                                                 --                .channel
			rf_sink_ready           => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                      --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	timer_1_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                      --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src6_ready,                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src6_valid,                                                   --                .valid
			cp_data                 => cmd_xbar_demux_001_src6_data,                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src6_startofpacket,                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src6_endofpacket,                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src6_channel,                                                 --                .channel
			rf_sink_ready           => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                      --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	pio_in_sw_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                        --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                    --       clk_reset.reset
			m0_address              => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src7_ready,                                                     --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src7_valid,                                                     --                .valid
			cp_data                 => cmd_xbar_demux_001_src7_data,                                                      --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src7_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src7_endofpacket,                                               --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src7_channel,                                                   --                .channel
			rf_sink_ready           => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                              --     (terminated)
			m0_writeresponserequest => open,                                                                              --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                --     (terminated)
		);

	pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                        --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                    -- clk_reset.reset
			in_data           => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                              -- (terminated)
			csr_read          => '0',                                                                               -- (terminated)
			csr_write         => '0',                                                                               -- (terminated)
			csr_readdata      => open,                                                                              -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                -- (terminated)
			almost_full_data  => open,                                                                              -- (terminated)
			almost_empty_data => open,                                                                              -- (terminated)
			in_empty          => '0',                                                                               -- (terminated)
			out_empty         => open,                                                                              -- (terminated)
			in_error          => '0',                                                                               -- (terminated)
			out_error         => open,                                                                              -- (terminated)
			in_channel        => '0',                                                                               -- (terminated)
			out_channel       => open                                                                               -- (terminated)
		);

	pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                              --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                          --       clk_reset.reset
			m0_address              => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src8_ready,                                                           --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src8_valid,                                                           --                .valid
			cp_data                 => cmd_xbar_demux_001_src8_data,                                                            --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src8_startofpacket,                                                   --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src8_endofpacket,                                                     --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src8_channel,                                                         --                .channel
			rf_sink_ready           => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                    --     (terminated)
			m0_writeresponserequest => open,                                                                                    --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                      --     (terminated)
		);

	pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                              --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                          -- clk_reset.reset
			in_data           => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                    -- (terminated)
			csr_read          => '0',                                                                                     -- (terminated)
			csr_write         => '0',                                                                                     -- (terminated)
			csr_readdata      => open,                                                                                    -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                      -- (terminated)
			almost_full_data  => open,                                                                                    -- (terminated)
			almost_empty_data => open,                                                                                    -- (terminated)
			in_empty          => '0',                                                                                     -- (terminated)
			out_empty         => open,                                                                                    -- (terminated)
			in_error          => '0',                                                                                     -- (terminated)
			out_error         => open,                                                                                    -- (terminated)
			in_channel        => '0',                                                                                     -- (terminated)
			out_channel       => open                                                                                     -- (terminated)
		);

	pio_in_ext_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                     --       clk_reset.reset
			m0_address              => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src9_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src9_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_demux_001_src9_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src9_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src9_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src9_channel,                                                    --                .channel
			rf_sink_ready           => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                 --     (terminated)
		);

	pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			in_data           => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                               -- (terminated)
			csr_read          => '0',                                                                                -- (terminated)
			csr_write         => '0',                                                                                -- (terminated)
			csr_readdata      => open,                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                 -- (terminated)
			almost_full_data  => open,                                                                               -- (terminated)
			almost_empty_data => open,                                                                               -- (terminated)
			in_empty          => '0',                                                                                -- (terminated)
			out_empty         => open,                                                                               -- (terminated)
			in_error          => '0',                                                                                -- (terminated)
			out_error         => open,                                                                               -- (terminated)
			in_channel        => '0',                                                                                -- (terminated)
			out_channel       => open                                                                                -- (terminated)
		);

	pio_out_red_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                          --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                      --       clk_reset.reset
			m0_address              => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_out_red_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src10_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src10_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_demux_001_src10_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src10_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src10_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src10_channel,                                                    --                .channel
			rf_sink_ready           => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                --     (terminated)
			m0_writeresponserequest => open,                                                                                --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                  --     (terminated)
		);

	pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                          --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                      -- clk_reset.reset
			in_data           => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                -- (terminated)
			csr_read          => '0',                                                                                 -- (terminated)
			csr_write         => '0',                                                                                 -- (terminated)
			csr_readdata      => open,                                                                                -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                  -- (terminated)
			almost_full_data  => open,                                                                                -- (terminated)
			almost_empty_data => open,                                                                                -- (terminated)
			in_empty          => '0',                                                                                 -- (terminated)
			out_empty         => open,                                                                                -- (terminated)
			in_error          => '0',                                                                                 -- (terminated)
			out_error         => open,                                                                                -- (terminated)
			in_channel        => '0',                                                                                 -- (terminated)
			out_channel       => open                                                                                 -- (terminated)
		);

	pio_out_green_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                        --       clk_reset.reset
			m0_address              => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_out_green_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src11_ready,                                                        --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src11_valid,                                                        --                .valid
			cp_data                 => cmd_xbar_demux_001_src11_data,                                                         --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src11_startofpacket,                                                --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src11_endofpacket,                                                  --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src11_channel,                                                      --                .channel
			rf_sink_ready           => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                  --     (terminated)
			m0_writeresponserequest => open,                                                                                  --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                    --     (terminated)
		);

	pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			in_data           => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                  -- (terminated)
			csr_read          => '0',                                                                                   -- (terminated)
			csr_write         => '0',                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                    -- (terminated)
			almost_full_data  => open,                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                  -- (terminated)
			in_empty          => '0',                                                                                   -- (terminated)
			out_empty         => open,                                                                                  -- (terminated)
			in_error          => '0',                                                                                   -- (terminated)
			out_error         => open,                                                                                  -- (terminated)
			in_channel        => '0',                                                                                   -- (terminated)
			out_channel       => open                                                                                   -- (terminated)
		);

	pio_out_ext_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                          --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                      --       clk_reset.reset
			m0_address              => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src12_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src12_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_demux_001_src12_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src12_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src12_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src12_channel,                                                    --                .channel
			rf_sink_ready           => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                --     (terminated)
			m0_writeresponserequest => open,                                                                                --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                  --     (terminated)
		);

	pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                          --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                      -- clk_reset.reset
			in_data           => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                -- (terminated)
			csr_read          => '0',                                                                                 -- (terminated)
			csr_write         => '0',                                                                                 -- (terminated)
			csr_readdata      => open,                                                                                -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                  -- (terminated)
			almost_full_data  => open,                                                                                -- (terminated)
			almost_empty_data => open,                                                                                -- (terminated)
			in_empty          => '0',                                                                                 -- (terminated)
			out_empty         => open,                                                                                -- (terminated)
			in_error          => '0',                                                                                 -- (terminated)
			out_error         => open,                                                                                -- (terminated)
			in_channel        => '0',                                                                                 -- (terminated)
			out_channel       => open                                                                                 -- (terminated)
		);

	pio_async_reset_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                              --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                          --       clk_reset.reset
			m0_address              => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src13_ready,                                                          --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src13_valid,                                                          --                .valid
			cp_data                 => cmd_xbar_demux_001_src13_data,                                                           --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src13_startofpacket,                                                  --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src13_endofpacket,                                                    --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src13_channel,                                                        --                .channel
			rf_sink_ready           => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                    --     (terminated)
			m0_writeresponserequest => open,                                                                                    --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                      --     (terminated)
		);

	pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                              --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                          -- clk_reset.reset
			in_data           => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                    -- (terminated)
			csr_read          => '0',                                                                                     -- (terminated)
			csr_write         => '0',                                                                                     -- (terminated)
			csr_readdata      => open,                                                                                    -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                      -- (terminated)
			almost_full_data  => open,                                                                                    -- (terminated)
			almost_empty_data => open,                                                                                    -- (terminated)
			in_empty          => '0',                                                                                     -- (terminated)
			out_empty         => open,                                                                                    -- (terminated)
			in_error          => '0',                                                                                     -- (terminated)
			out_error         => open,                                                                                    -- (terminated)
			in_channel        => '0',                                                                                     -- (terminated)
			out_channel       => open                                                                                     -- (terminated)
		);

	pio_en_mux_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                     --       clk_reset.reset
			m0_address              => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src14_ready,                                                     --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src14_valid,                                                     --                .valid
			cp_data                 => cmd_xbar_demux_001_src14_data,                                                      --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src14_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src14_endofpacket,                                               --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src14_channel,                                                   --                .channel
			rf_sink_ready           => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                 --     (terminated)
		);

	pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			in_data           => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                               -- (terminated)
			csr_read          => '0',                                                                                -- (terminated)
			csr_write         => '0',                                                                                -- (terminated)
			csr_readdata      => open,                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                 -- (terminated)
			almost_full_data  => open,                                                                               -- (terminated)
			almost_empty_data => open,                                                                               -- (terminated)
			in_empty          => '0',                                                                                -- (terminated)
			out_empty         => open,                                                                               -- (terminated)
			in_error          => '0',                                                                                -- (terminated)
			out_error         => open,                                                                               -- (terminated)
			in_channel        => '0',                                                                                -- (terminated)
			out_channel       => open                                                                                -- (terminated)
		);

	pio_direc_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                        --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                    --       clk_reset.reset
			m0_address              => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_direc_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_direc_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_direc_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_direc_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_direc_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_direc_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src15_ready,                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src15_valid,                                                    --                .valid
			cp_data                 => cmd_xbar_demux_001_src15_data,                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src15_startofpacket,                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src15_endofpacket,                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src15_channel,                                                  --                .channel
			rf_sink_ready           => pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_direc_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_direc_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_direc_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_direc_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_direc_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_direc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_direc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_direc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_direc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_direc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_direc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                              --     (terminated)
			m0_writeresponserequest => open,                                                                              --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                --     (terminated)
		);

	pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                        --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                    -- clk_reset.reset
			in_data           => pio_direc_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_direc_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_direc_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_direc_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_direc_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_direc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                              -- (terminated)
			csr_read          => '0',                                                                               -- (terminated)
			csr_write         => '0',                                                                               -- (terminated)
			csr_readdata      => open,                                                                              -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                -- (terminated)
			almost_full_data  => open,                                                                              -- (terminated)
			almost_empty_data => open,                                                                              -- (terminated)
			in_empty          => '0',                                                                               -- (terminated)
			out_empty         => open,                                                                              -- (terminated)
			in_error          => '0',                                                                               -- (terminated)
			out_error         => open,                                                                              -- (terminated)
			in_channel        => '0',                                                                               -- (terminated)
			out_channel       => open                                                                               -- (terminated)
		);

	pio_direc_ram_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                        --       clk_reset.reset
			m0_address              => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src16_ready,                                                        --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src16_valid,                                                        --                .valid
			cp_data                 => cmd_xbar_demux_001_src16_data,                                                         --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src16_startofpacket,                                                --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src16_endofpacket,                                                  --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src16_channel,                                                      --                .channel
			rf_sink_ready           => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                  --     (terminated)
			m0_writeresponserequest => open,                                                                                  --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                    --     (terminated)
		);

	pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			in_data           => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                  -- (terminated)
			csr_read          => '0',                                                                                   -- (terminated)
			csr_write         => '0',                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                    -- (terminated)
			almost_full_data  => open,                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                  -- (terminated)
			in_empty          => '0',                                                                                   -- (terminated)
			out_empty         => open,                                                                                  -- (terminated)
			in_error          => '0',                                                                                   -- (terminated)
			out_error         => open,                                                                                  -- (terminated)
			in_channel        => '0',                                                                                   -- (terminated)
			out_channel       => open                                                                                   -- (terminated)
		);

	pio_wr_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                     --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                 --       clk_reset.reset
			m0_address              => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_wr_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_wr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_wr_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_wr_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_wr_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_wr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src17_ready,                                                 --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src17_valid,                                                 --                .valid
			cp_data                 => cmd_xbar_demux_001_src17_data,                                                  --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src17_startofpacket,                                         --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src17_endofpacket,                                           --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src17_channel,                                               --                .channel
			rf_sink_ready           => pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_wr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_wr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_wr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_wr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_wr_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_wr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_wr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_wr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_wr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_wr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_wr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                             --     (terminated)
		);

	pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                     --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			in_data           => pio_wr_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_wr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_wr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_wr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_wr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_wr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                           -- (terminated)
			csr_read          => '0',                                                                            -- (terminated)
			csr_write         => '0',                                                                            -- (terminated)
			csr_readdata      => open,                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                             -- (terminated)
			almost_full_data  => open,                                                                           -- (terminated)
			almost_empty_data => open,                                                                           -- (terminated)
			in_empty          => '0',                                                                            -- (terminated)
			out_empty         => open,                                                                           -- (terminated)
			in_error          => '0',                                                                            -- (terminated)
			out_error         => open,                                                                           -- (terminated)
			in_channel        => '0',                                                                            -- (terminated)
			out_channel       => open                                                                            -- (terminated)
		);

	pio_sel_salida_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                             --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                         --       clk_reset.reset
			m0_address              => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src18_ready,                                                         --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src18_valid,                                                         --                .valid
			cp_data                 => cmd_xbar_demux_001_src18_data,                                                          --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src18_startofpacket,                                                 --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src18_endofpacket,                                                   --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src18_channel,                                                       --                .channel
			rf_sink_ready           => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                   --     (terminated)
			m0_writeresponserequest => open,                                                                                   --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                     --     (terminated)
		);

	pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                             --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                         -- clk_reset.reset
			in_data           => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                   -- (terminated)
			csr_read          => '0',                                                                                    -- (terminated)
			csr_write         => '0',                                                                                    -- (terminated)
			csr_readdata      => open,                                                                                   -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                     -- (terminated)
			almost_full_data  => open,                                                                                   -- (terminated)
			almost_empty_data => open,                                                                                   -- (terminated)
			in_empty          => '0',                                                                                    -- (terminated)
			out_empty         => open,                                                                                   -- (terminated)
			in_error          => '0',                                                                                    -- (terminated)
			out_error         => open,                                                                                   -- (terminated)
			in_channel        => '0',                                                                                    -- (terminated)
			out_channel       => open                                                                                    -- (terminated)
		);

	pio_datos_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                        --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                    --       clk_reset.reset
			m0_address              => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_datos_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_datos_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_datos_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_datos_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_datos_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_datos_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src19_ready,                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src19_valid,                                                    --                .valid
			cp_data                 => cmd_xbar_demux_001_src19_data,                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src19_startofpacket,                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src19_endofpacket,                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src19_channel,                                                  --                .channel
			rf_sink_ready           => pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_datos_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_datos_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_datos_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_datos_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_datos_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_datos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_datos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_datos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_datos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_datos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_datos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                              --     (terminated)
			m0_writeresponserequest => open,                                                                              --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                --     (terminated)
		);

	pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                        --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                    -- clk_reset.reset
			in_data           => pio_datos_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_datos_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_datos_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_datos_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_datos_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_datos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                              -- (terminated)
			csr_read          => '0',                                                                               -- (terminated)
			csr_write         => '0',                                                                               -- (terminated)
			csr_readdata      => open,                                                                              -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                -- (terminated)
			almost_full_data  => open,                                                                              -- (terminated)
			almost_empty_data => open,                                                                              -- (terminated)
			in_empty          => '0',                                                                               -- (terminated)
			out_empty         => open,                                                                              -- (terminated)
			in_error          => '0',                                                                               -- (terminated)
			out_error         => open,                                                                              -- (terminated)
			in_channel        => '0',                                                                               -- (terminated)
			out_channel       => open                                                                               -- (terminated)
		);

	pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                                --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                            --       clk_reset.reset
			m0_address              => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src20_ready,                                                            --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src20_valid,                                                            --                .valid
			cp_data                 => cmd_xbar_demux_001_src20_data,                                                             --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src20_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src20_endofpacket,                                                      --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src20_channel,                                                          --                .channel
			rf_sink_ready           => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                      --     (terminated)
			m0_writeresponserequest => open,                                                                                      --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                        --     (terminated)
		);

	pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                                --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			in_data           => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                      -- (terminated)
			csr_read          => '0',                                                                                       -- (terminated)
			csr_write         => '0',                                                                                       -- (terminated)
			csr_readdata      => open,                                                                                      -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                        -- (terminated)
			almost_full_data  => open,                                                                                      -- (terminated)
			almost_empty_data => open,                                                                                      -- (terminated)
			in_empty          => '0',                                                                                       -- (terminated)
			out_empty         => open,                                                                                      -- (terminated)
			in_error          => '0',                                                                                       -- (terminated)
			out_error         => open,                                                                                      -- (terminated)
			in_channel        => '0',                                                                                       -- (terminated)
			out_channel       => open                                                                                       -- (terminated)
		);

	pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                                --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                            --       clk_reset.reset
			m0_address              => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src21_ready,                                                            --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src21_valid,                                                            --                .valid
			cp_data                 => cmd_xbar_demux_001_src21_data,                                                             --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src21_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src21_endofpacket,                                                      --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src21_channel,                                                          --                .channel
			rf_sink_ready           => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                      --     (terminated)
			m0_writeresponserequest => open,                                                                                      --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                        --     (terminated)
		);

	pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                                --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			in_data           => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                      -- (terminated)
			csr_read          => '0',                                                                                       -- (terminated)
			csr_write         => '0',                                                                                       -- (terminated)
			csr_readdata      => open,                                                                                      -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                        -- (terminated)
			almost_full_data  => open,                                                                                      -- (terminated)
			almost_empty_data => open,                                                                                      -- (terminated)
			in_empty          => '0',                                                                                       -- (terminated)
			out_empty         => open,                                                                                      -- (terminated)
			in_error          => '0',                                                                                       -- (terminated)
			out_error         => open,                                                                                      -- (terminated)
			in_channel        => '0',                                                                                       -- (terminated)
			out_channel       => open                                                                                       -- (terminated)
		);

	pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                                --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                            --       clk_reset.reset
			m0_address              => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src22_ready,                                                            --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src22_valid,                                                            --                .valid
			cp_data                 => cmd_xbar_demux_001_src22_data,                                                             --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src22_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src22_endofpacket,                                                      --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src22_channel,                                                          --                .channel
			rf_sink_ready           => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                      --     (terminated)
			m0_writeresponserequest => open,                                                                                      --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                        --     (terminated)
		);

	pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                                --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			in_data           => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                      -- (terminated)
			csr_read          => '0',                                                                                       -- (terminated)
			csr_write         => '0',                                                                                       -- (terminated)
			csr_readdata      => open,                                                                                      -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                        -- (terminated)
			almost_full_data  => open,                                                                                      -- (terminated)
			almost_empty_data => open,                                                                                      -- (terminated)
			in_empty          => '0',                                                                                       -- (terminated)
			out_empty         => open,                                                                                      -- (terminated)
			in_error          => '0',                                                                                       -- (terminated)
			out_error         => open,                                                                                      -- (terminated)
			in_channel        => '0',                                                                                       -- (terminated)
			out_channel       => open                                                                                       -- (terminated)
		);

	pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                                --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                            --       clk_reset.reset
			m0_address              => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src23_ready,                                                            --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src23_valid,                                                            --                .valid
			cp_data                 => cmd_xbar_demux_001_src23_data,                                                             --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src23_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src23_endofpacket,                                                      --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src23_channel,                                                          --                .channel
			rf_sink_ready           => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                      --     (terminated)
			m0_writeresponserequest => open,                                                                                      --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                        --     (terminated)
		);

	pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                                --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			in_data           => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                      -- (terminated)
			csr_read          => '0',                                                                                       -- (terminated)
			csr_write         => '0',                                                                                       -- (terminated)
			csr_readdata      => open,                                                                                      -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                        -- (terminated)
			almost_full_data  => open,                                                                                      -- (terminated)
			almost_empty_data => open,                                                                                      -- (terminated)
			in_empty          => '0',                                                                                       -- (terminated)
			out_empty         => open,                                                                                      -- (terminated)
			in_error          => '0',                                                                                       -- (terminated)
			out_error         => open,                                                                                      -- (terminated)
			in_channel        => '0',                                                                                       -- (terminated)
			out_channel       => open                                                                                       -- (terminated)
		);

	pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                                --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                            --       clk_reset.reset
			m0_address              => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src24_ready,                                                            --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src24_valid,                                                            --                .valid
			cp_data                 => cmd_xbar_demux_001_src24_data,                                                             --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src24_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src24_endofpacket,                                                      --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src24_channel,                                                          --                .channel
			rf_sink_ready           => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                      --     (terminated)
			m0_writeresponserequest => open,                                                                                      --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                        --     (terminated)
		);

	pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                                --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			in_data           => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                      -- (terminated)
			csr_read          => '0',                                                                                       -- (terminated)
			csr_write         => '0',                                                                                       -- (terminated)
			csr_readdata      => open,                                                                                      -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                        -- (terminated)
			almost_full_data  => open,                                                                                      -- (terminated)
			almost_empty_data => open,                                                                                      -- (terminated)
			in_empty          => '0',                                                                                       -- (terminated)
			out_empty         => open,                                                                                      -- (terminated)
			in_error          => '0',                                                                                       -- (terminated)
			out_error         => open,                                                                                      -- (terminated)
			in_channel        => '0',                                                                                       -- (terminated)
			out_channel       => open                                                                                       -- (terminated)
		);

	pio_captura_0_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                        --       clk_reset.reset
			m0_address              => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src25_ready,                                                        --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src25_valid,                                                        --                .valid
			cp_data                 => cmd_xbar_demux_001_src25_data,                                                         --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src25_startofpacket,                                                --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src25_endofpacket,                                                  --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src25_channel,                                                      --                .channel
			rf_sink_ready           => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                  --     (terminated)
			m0_writeresponserequest => open,                                                                                  --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                    --     (terminated)
		);

	pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			in_data           => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                  -- (terminated)
			csr_read          => '0',                                                                                   -- (terminated)
			csr_write         => '0',                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                    -- (terminated)
			almost_full_data  => open,                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                  -- (terminated)
			in_empty          => '0',                                                                                   -- (terminated)
			out_empty         => open,                                                                                  -- (terminated)
			in_error          => '0',                                                                                   -- (terminated)
			out_error         => open,                                                                                  -- (terminated)
			in_channel        => '0',                                                                                   -- (terminated)
			out_channel       => open                                                                                   -- (terminated)
		);

	pio_captura_1_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                        --       clk_reset.reset
			m0_address              => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src26_ready,                                                        --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src26_valid,                                                        --                .valid
			cp_data                 => cmd_xbar_demux_001_src26_data,                                                         --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src26_startofpacket,                                                --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src26_endofpacket,                                                  --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src26_channel,                                                      --                .channel
			rf_sink_ready           => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                  --     (terminated)
			m0_writeresponserequest => open,                                                                                  --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                    --     (terminated)
		);

	pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			in_data           => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                  -- (terminated)
			csr_read          => '0',                                                                                   -- (terminated)
			csr_write         => '0',                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                    -- (terminated)
			almost_full_data  => open,                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                  -- (terminated)
			in_empty          => '0',                                                                                   -- (terminated)
			out_empty         => open,                                                                                  -- (terminated)
			in_error          => '0',                                                                                   -- (terminated)
			out_error         => open,                                                                                  -- (terminated)
			in_channel        => '0',                                                                                   -- (terminated)
			out_channel       => open                                                                                   -- (terminated)
		);

	pio_captura_2_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                        --       clk_reset.reset
			m0_address              => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src27_ready,                                                        --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src27_valid,                                                        --                .valid
			cp_data                 => cmd_xbar_demux_001_src27_data,                                                         --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src27_startofpacket,                                                --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src27_endofpacket,                                                  --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src27_channel,                                                      --                .channel
			rf_sink_ready           => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                  --     (terminated)
			m0_writeresponserequest => open,                                                                                  --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                    --     (terminated)
		);

	pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			in_data           => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                  -- (terminated)
			csr_read          => '0',                                                                                   -- (terminated)
			csr_write         => '0',                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                    -- (terminated)
			almost_full_data  => open,                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                  -- (terminated)
			in_empty          => '0',                                                                                   -- (terminated)
			out_empty         => open,                                                                                  -- (terminated)
			in_error          => '0',                                                                                   -- (terminated)
			out_error         => open,                                                                                  -- (terminated)
			in_channel        => '0',                                                                                   -- (terminated)
			out_channel       => open                                                                                   -- (terminated)
		);

	pio_captura_3_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                        --       clk_reset.reset
			m0_address              => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src28_ready,                                                        --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src28_valid,                                                        --                .valid
			cp_data                 => cmd_xbar_demux_001_src28_data,                                                         --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src28_startofpacket,                                                --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src28_endofpacket,                                                  --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src28_channel,                                                      --                .channel
			rf_sink_ready           => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                  --     (terminated)
			m0_writeresponserequest => open,                                                                                  --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                    --     (terminated)
		);

	pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			in_data           => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                  -- (terminated)
			csr_read          => '0',                                                                                   -- (terminated)
			csr_write         => '0',                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                    -- (terminated)
			almost_full_data  => open,                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                  -- (terminated)
			in_empty          => '0',                                                                                   -- (terminated)
			out_empty         => open,                                                                                  -- (terminated)
			in_error          => '0',                                                                                   -- (terminated)
			out_error         => open,                                                                                  -- (terminated)
			in_channel        => '0',                                                                                   -- (terminated)
			out_channel       => open                                                                                   -- (terminated)
		);

	pio_captura_4_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                        --       clk_reset.reset
			m0_address              => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src29_ready,                                                        --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src29_valid,                                                        --                .valid
			cp_data                 => cmd_xbar_demux_001_src29_data,                                                         --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src29_startofpacket,                                                --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src29_endofpacket,                                                  --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src29_channel,                                                      --                .channel
			rf_sink_ready           => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                  --     (terminated)
			m0_writeresponserequest => open,                                                                                  --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                    --     (terminated)
		);

	pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			in_data           => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                  -- (terminated)
			csr_read          => '0',                                                                                   -- (terminated)
			csr_write         => '0',                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                    -- (terminated)
			almost_full_data  => open,                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                  -- (terminated)
			in_empty          => '0',                                                                                   -- (terminated)
			out_empty         => open,                                                                                  -- (terminated)
			in_error          => '0',                                                                                   -- (terminated)
			out_error         => open,                                                                                  -- (terminated)
			in_channel        => '0',                                                                                   -- (terminated)
			out_channel       => open                                                                                   -- (terminated)
		);

	pio_in_32_s1_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                        --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                    --       clk_reset.reset
			m0_address              => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_in_32_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src30_ready,                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src30_valid,                                                    --                .valid
			cp_data                 => cmd_xbar_demux_001_src30_data,                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src30_startofpacket,                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src30_endofpacket,                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src30_channel,                                                  --                .channel
			rf_sink_ready           => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                              --     (terminated)
			m0_writeresponserequest => open,                                                                              --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                --     (terminated)
		);

	pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                        --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                    -- clk_reset.reset
			in_data           => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                              -- (terminated)
			csr_read          => '0',                                                                               -- (terminated)
			csr_write         => '0',                                                                               -- (terminated)
			csr_readdata      => open,                                                                              -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                -- (terminated)
			almost_full_data  => open,                                                                              -- (terminated)
			almost_empty_data => open,                                                                              -- (terminated)
			in_empty          => '0',                                                                               -- (terminated)
			out_empty         => open,                                                                              -- (terminated)
			in_error          => '0',                                                                               -- (terminated)
			out_error         => open,                                                                              -- (terminated)
			in_channel        => '0',                                                                               -- (terminated)
			out_channel       => open                                                                               -- (terminated)
		);

	lcd_control_slave_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                             --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                         --       clk_reset.reset
			m0_address              => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src31_ready,                                                         --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src31_valid,                                                         --                .valid
			cp_data                 => cmd_xbar_demux_001_src31_data,                                                          --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src31_startofpacket,                                                 --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src31_endofpacket,                                                   --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src31_channel,                                                       --                .channel
			rf_sink_ready           => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                   --     (terminated)
			m0_writeresponserequest => open,                                                                                   --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                     --     (terminated)
		);

	lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                             --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                         -- clk_reset.reset
			in_data           => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                   -- (terminated)
			csr_read          => '0',                                                                                    -- (terminated)
			csr_write         => '0',                                                                                    -- (terminated)
			csr_readdata      => open,                                                                                   -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                     -- (terminated)
			almost_full_data  => open,                                                                                   -- (terminated)
			almost_empty_data => open,                                                                                   -- (terminated)
			in_empty          => '0',                                                                                    -- (terminated)
			out_empty         => open,                                                                                   -- (terminated)
			in_error          => '0',                                                                                    -- (terminated)
			out_error         => open,                                                                                   -- (terminated)
			in_channel        => '0',                                                                                    -- (terminated)
			out_channel       => open                                                                                    -- (terminated)
		);

	dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 97,
			PKT_PROTECTION_L          => 95,
			PKT_RESPONSE_STATUS_H     => 103,
			PKT_RESPONSE_STATUS_L     => 102,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 33,
			ST_DATA_W                 => 104,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => pll_c0_clk,                                                                                  --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                              --       clk_reset.reset
			m0_address              => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src32_ready,                                                              --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src32_valid,                                                              --                .valid
			cp_data                 => cmd_xbar_demux_001_src32_data,                                                               --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src32_startofpacket,                                                      --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src32_endofpacket,                                                        --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src32_channel,                                                            --                .channel
			rf_sink_ready           => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                          --     (terminated)
		);

	dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component niosiimicro_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 105,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => pll_c0_clk,                                                                                  --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                              -- clk_reset.reset
			in_data           => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                        -- (terminated)
			csr_read          => '0',                                                                                         -- (terminated)
			csr_write         => '0',                                                                                         -- (terminated)
			csr_readdata      => open,                                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                          -- (terminated)
			almost_full_data  => open,                                                                                        -- (terminated)
			almost_empty_data => open,                                                                                        -- (terminated)
			in_empty          => '0',                                                                                         -- (terminated)
			out_empty         => open,                                                                                        -- (terminated)
			in_error          => '0',                                                                                         -- (terminated)
			out_error         => open,                                                                                        -- (terminated)
			in_channel        => '0',                                                                                         -- (terminated)
			out_channel       => open                                                                                         -- (terminated)
		);

	addr_router : component NIOSIImicro_addr_router
		port map (
			sink_ready         => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                         --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                              --       src.ready
			src_valid          => addr_router_src_valid,                                                              --          .valid
			src_data           => addr_router_src_data,                                                               --          .data
			src_channel        => addr_router_src_channel,                                                            --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                         --          .endofpacket
		);

	addr_router_001 : component NIOSIImicro_addr_router_001
		port map (
			sink_ready         => cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                   --       src.ready
			src_valid          => addr_router_001_src_valid,                                                   --          .valid
			src_data           => addr_router_001_src_data,                                                    --          .data
			src_channel        => addr_router_001_src_channel,                                                 --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                           --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                              --          .endofpacket
		);

	id_router : component NIOSIImicro_id_router
		port map (
			sink_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                       --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                              --       src.ready
			src_valid          => id_router_src_valid,                                                              --          .valid
			src_data           => id_router_src_data,                                                               --          .data
			src_channel        => id_router_src_channel,                                                            --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                         --          .endofpacket
		);

	id_router_001 : component NIOSIImicro_id_router_001
		port map (
			sink_ready         => sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sdram_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                          --       clk.clk
			reset              => rst_controller_reset_out_reset,                                      -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                             --       src.ready
			src_valid          => id_router_001_src_valid,                                             --          .valid
			src_data           => id_router_001_src_data,                                              --          .data
			src_channel        => id_router_001_src_channel,                                           --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                     --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                        --          .endofpacket
		);

	id_router_002 : component NIOSIImicro_id_router
		port map (
			sink_ready         => system_id_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => system_id_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => system_id_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => system_id_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => system_id_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                         --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                                            --       src.ready
			src_valid          => id_router_002_src_valid,                                                            --          .valid
			src_data           => id_router_002_src_data,                                                             --          .data
			src_channel        => id_router_002_src_channel,                                                          --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                                    --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                                       --          .endofpacket
		);

	id_router_003 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50_clk,                                                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                       -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                  --       src.ready
			src_valid          => id_router_003_src_valid,                                                  --          .valid
			src_data           => id_router_003_src_data,                                                   --          .data
			src_channel        => id_router_003_src_channel,                                                --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                          --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                             --          .endofpacket
		);

	id_router_004 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                        --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                    -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                                           --       src.ready
			src_valid          => id_router_004_src_valid,                                                           --          .valid
			src_data           => id_router_004_src_data,                                                            --          .data
			src_channel        => id_router_004_src_channel,                                                         --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                                   --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                                      --          .endofpacket
		);

	id_router_005 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                               --       src.ready
			src_valid          => id_router_005_src_valid,                                               --          .valid
			src_data           => id_router_005_src_data,                                                --          .data
			src_channel        => id_router_005_src_channel,                                             --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                          --          .endofpacket
		);

	id_router_006 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                               --       src.ready
			src_valid          => id_router_006_src_valid,                                               --          .valid
			src_data           => id_router_006_src_data,                                                --          .data
			src_channel        => id_router_006_src_channel,                                             --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                          --          .endofpacket
		);

	id_router_007 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_in_sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                          -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                                 --       src.ready
			src_valid          => id_router_007_src_valid,                                                 --          .valid
			src_data           => id_router_007_src_data,                                                  --          .data
			src_channel        => id_router_007_src_channel,                                               --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                         --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                            --          .endofpacket
		);

	id_router_008 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_in_key_edge_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                    --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                -- clk_reset.reset
			src_ready          => id_router_008_src_ready,                                                       --       src.ready
			src_valid          => id_router_008_src_valid,                                                       --          .valid
			src_data           => id_router_008_src_data,                                                        --          .data
			src_channel        => id_router_008_src_channel,                                                     --          .channel
			src_startofpacket  => id_router_008_src_startofpacket,                                               --          .startofpacket
			src_endofpacket    => id_router_008_src_endofpacket                                                  --          .endofpacket
		);

	id_router_009 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_in_ext_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                           -- clk_reset.reset
			src_ready          => id_router_009_src_ready,                                                  --       src.ready
			src_valid          => id_router_009_src_valid,                                                  --          .valid
			src_data           => id_router_009_src_data,                                                   --          .data
			src_channel        => id_router_009_src_channel,                                                --          .channel
			src_startofpacket  => id_router_009_src_startofpacket,                                          --          .startofpacket
			src_endofpacket    => id_router_009_src_endofpacket                                             --          .endofpacket
		);

	id_router_010 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_out_red_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                --       clk.clk
			reset              => rst_controller_reset_out_reset,                                            -- clk_reset.reset
			src_ready          => id_router_010_src_ready,                                                   --       src.ready
			src_valid          => id_router_010_src_valid,                                                   --          .valid
			src_data           => id_router_010_src_data,                                                    --          .data
			src_channel        => id_router_010_src_channel,                                                 --          .channel
			src_startofpacket  => id_router_010_src_startofpacket,                                           --          .startofpacket
			src_endofpacket    => id_router_010_src_endofpacket                                              --          .endofpacket
		);

	id_router_011 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_out_green_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => id_router_011_src_ready,                                                     --       src.ready
			src_valid          => id_router_011_src_valid,                                                     --          .valid
			src_data           => id_router_011_src_data,                                                      --          .data
			src_channel        => id_router_011_src_channel,                                                   --          .channel
			src_startofpacket  => id_router_011_src_startofpacket,                                             --          .startofpacket
			src_endofpacket    => id_router_011_src_endofpacket                                                --          .endofpacket
		);

	id_router_012 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_out_ext_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                --       clk.clk
			reset              => rst_controller_reset_out_reset,                                            -- clk_reset.reset
			src_ready          => id_router_012_src_ready,                                                   --       src.ready
			src_valid          => id_router_012_src_valid,                                                   --          .valid
			src_data           => id_router_012_src_data,                                                    --          .data
			src_channel        => id_router_012_src_channel,                                                 --          .channel
			src_startofpacket  => id_router_012_src_startofpacket,                                           --          .startofpacket
			src_endofpacket    => id_router_012_src_endofpacket                                              --          .endofpacket
		);

	id_router_013 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_async_reset_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                    --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                -- clk_reset.reset
			src_ready          => id_router_013_src_ready,                                                       --       src.ready
			src_valid          => id_router_013_src_valid,                                                       --          .valid
			src_data           => id_router_013_src_data,                                                        --          .data
			src_channel        => id_router_013_src_channel,                                                     --          .channel
			src_startofpacket  => id_router_013_src_startofpacket,                                               --          .startofpacket
			src_endofpacket    => id_router_013_src_endofpacket                                                  --          .endofpacket
		);

	id_router_014 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_en_mux_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                           -- clk_reset.reset
			src_ready          => id_router_014_src_ready,                                                  --       src.ready
			src_valid          => id_router_014_src_valid,                                                  --          .valid
			src_data           => id_router_014_src_data,                                                   --          .data
			src_channel        => id_router_014_src_channel,                                                --          .channel
			src_startofpacket  => id_router_014_src_startofpacket,                                          --          .startofpacket
			src_endofpacket    => id_router_014_src_endofpacket                                             --          .endofpacket
		);

	id_router_015 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_direc_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_direc_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_direc_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_direc_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_direc_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                          -- clk_reset.reset
			src_ready          => id_router_015_src_ready,                                                 --       src.ready
			src_valid          => id_router_015_src_valid,                                                 --          .valid
			src_data           => id_router_015_src_data,                                                  --          .data
			src_channel        => id_router_015_src_channel,                                               --          .channel
			src_startofpacket  => id_router_015_src_startofpacket,                                         --          .startofpacket
			src_endofpacket    => id_router_015_src_endofpacket                                            --          .endofpacket
		);

	id_router_016 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_direc_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => id_router_016_src_ready,                                                     --       src.ready
			src_valid          => id_router_016_src_valid,                                                     --          .valid
			src_data           => id_router_016_src_data,                                                      --          .data
			src_channel        => id_router_016_src_channel,                                                   --          .channel
			src_startofpacket  => id_router_016_src_startofpacket,                                             --          .startofpacket
			src_endofpacket    => id_router_016_src_endofpacket                                                --          .endofpacket
		);

	id_router_017 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_wr_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_wr_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_wr_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_wr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_wr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                           --       clk.clk
			reset              => rst_controller_reset_out_reset,                                       -- clk_reset.reset
			src_ready          => id_router_017_src_ready,                                              --       src.ready
			src_valid          => id_router_017_src_valid,                                              --          .valid
			src_data           => id_router_017_src_data,                                               --          .data
			src_channel        => id_router_017_src_channel,                                            --          .channel
			src_startofpacket  => id_router_017_src_startofpacket,                                      --          .startofpacket
			src_endofpacket    => id_router_017_src_endofpacket                                         --          .endofpacket
		);

	id_router_018 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_sel_salida_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                   --       clk.clk
			reset              => rst_controller_reset_out_reset,                                               -- clk_reset.reset
			src_ready          => id_router_018_src_ready,                                                      --       src.ready
			src_valid          => id_router_018_src_valid,                                                      --          .valid
			src_data           => id_router_018_src_data,                                                       --          .data
			src_channel        => id_router_018_src_channel,                                                    --          .channel
			src_startofpacket  => id_router_018_src_startofpacket,                                              --          .startofpacket
			src_endofpacket    => id_router_018_src_endofpacket                                                 --          .endofpacket
		);

	id_router_019 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_datos_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_datos_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_datos_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_datos_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_datos_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                          -- clk_reset.reset
			src_ready          => id_router_019_src_ready,                                                 --       src.ready
			src_valid          => id_router_019_src_valid,                                                 --          .valid
			src_data           => id_router_019_src_data,                                                  --          .data
			src_channel        => id_router_019_src_channel,                                               --          .channel
			src_startofpacket  => id_router_019_src_startofpacket,                                         --          .startofpacket
			src_endofpacket    => id_router_019_src_endofpacket                                            --          .endofpacket
		);

	id_router_020 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_compara_int_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                      --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			src_ready          => id_router_020_src_ready,                                                         --       src.ready
			src_valid          => id_router_020_src_valid,                                                         --          .valid
			src_data           => id_router_020_src_data,                                                          --          .data
			src_channel        => id_router_020_src_channel,                                                       --          .channel
			src_startofpacket  => id_router_020_src_startofpacket,                                                 --          .startofpacket
			src_endofpacket    => id_router_020_src_endofpacket                                                    --          .endofpacket
		);

	id_router_021 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_compara_int_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                      --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			src_ready          => id_router_021_src_ready,                                                         --       src.ready
			src_valid          => id_router_021_src_valid,                                                         --          .valid
			src_data           => id_router_021_src_data,                                                          --          .data
			src_channel        => id_router_021_src_channel,                                                       --          .channel
			src_startofpacket  => id_router_021_src_startofpacket,                                                 --          .startofpacket
			src_endofpacket    => id_router_021_src_endofpacket                                                    --          .endofpacket
		);

	id_router_022 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_compara_int_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                      --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			src_ready          => id_router_022_src_ready,                                                         --       src.ready
			src_valid          => id_router_022_src_valid,                                                         --          .valid
			src_data           => id_router_022_src_data,                                                          --          .data
			src_channel        => id_router_022_src_channel,                                                       --          .channel
			src_startofpacket  => id_router_022_src_startofpacket,                                                 --          .startofpacket
			src_endofpacket    => id_router_022_src_endofpacket                                                    --          .endofpacket
		);

	id_router_023 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_compara_int_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                      --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			src_ready          => id_router_023_src_ready,                                                         --       src.ready
			src_valid          => id_router_023_src_valid,                                                         --          .valid
			src_data           => id_router_023_src_data,                                                          --          .data
			src_channel        => id_router_023_src_channel,                                                       --          .channel
			src_startofpacket  => id_router_023_src_startofpacket,                                                 --          .startofpacket
			src_endofpacket    => id_router_023_src_endofpacket                                                    --          .endofpacket
		);

	id_router_024 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_compara_int_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                      --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			src_ready          => id_router_024_src_ready,                                                         --       src.ready
			src_valid          => id_router_024_src_valid,                                                         --          .valid
			src_data           => id_router_024_src_data,                                                          --          .data
			src_channel        => id_router_024_src_channel,                                                       --          .channel
			src_startofpacket  => id_router_024_src_startofpacket,                                                 --          .startofpacket
			src_endofpacket    => id_router_024_src_endofpacket                                                    --          .endofpacket
		);

	id_router_025 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_captura_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => id_router_025_src_ready,                                                     --       src.ready
			src_valid          => id_router_025_src_valid,                                                     --          .valid
			src_data           => id_router_025_src_data,                                                      --          .data
			src_channel        => id_router_025_src_channel,                                                   --          .channel
			src_startofpacket  => id_router_025_src_startofpacket,                                             --          .startofpacket
			src_endofpacket    => id_router_025_src_endofpacket                                                --          .endofpacket
		);

	id_router_026 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_captura_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => id_router_026_src_ready,                                                     --       src.ready
			src_valid          => id_router_026_src_valid,                                                     --          .valid
			src_data           => id_router_026_src_data,                                                      --          .data
			src_channel        => id_router_026_src_channel,                                                   --          .channel
			src_startofpacket  => id_router_026_src_startofpacket,                                             --          .startofpacket
			src_endofpacket    => id_router_026_src_endofpacket                                                --          .endofpacket
		);

	id_router_027 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_captura_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => id_router_027_src_ready,                                                     --       src.ready
			src_valid          => id_router_027_src_valid,                                                     --          .valid
			src_data           => id_router_027_src_data,                                                      --          .data
			src_channel        => id_router_027_src_channel,                                                   --          .channel
			src_startofpacket  => id_router_027_src_startofpacket,                                             --          .startofpacket
			src_endofpacket    => id_router_027_src_endofpacket                                                --          .endofpacket
		);

	id_router_028 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_captura_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => id_router_028_src_ready,                                                     --       src.ready
			src_valid          => id_router_028_src_valid,                                                     --          .valid
			src_data           => id_router_028_src_data,                                                      --          .data
			src_channel        => id_router_028_src_channel,                                                   --          .channel
			src_startofpacket  => id_router_028_src_startofpacket,                                             --          .startofpacket
			src_endofpacket    => id_router_028_src_endofpacket                                                --          .endofpacket
		);

	id_router_029 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_captura_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => id_router_029_src_ready,                                                     --       src.ready
			src_valid          => id_router_029_src_valid,                                                     --          .valid
			src_data           => id_router_029_src_data,                                                      --          .data
			src_channel        => id_router_029_src_channel,                                                   --          .channel
			src_startofpacket  => id_router_029_src_startofpacket,                                             --          .startofpacket
			src_endofpacket    => id_router_029_src_endofpacket                                                --          .endofpacket
		);

	id_router_030 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_in_32_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                          -- clk_reset.reset
			src_ready          => id_router_030_src_ready,                                                 --       src.ready
			src_valid          => id_router_030_src_valid,                                                 --          .valid
			src_data           => id_router_030_src_data,                                                  --          .data
			src_channel        => id_router_030_src_channel,                                               --          .channel
			src_startofpacket  => id_router_030_src_startofpacket,                                         --          .startofpacket
			src_endofpacket    => id_router_030_src_endofpacket                                            --          .endofpacket
		);

	id_router_031 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                   --       clk.clk
			reset              => rst_controller_reset_out_reset,                                               -- clk_reset.reset
			src_ready          => id_router_031_src_ready,                                                      --       src.ready
			src_valid          => id_router_031_src_valid,                                                      --          .valid
			src_data           => id_router_031_src_data,                                                       --          .data
			src_channel        => id_router_031_src_channel,                                                    --          .channel
			src_startofpacket  => id_router_031_src_startofpacket,                                              --          .startofpacket
			src_endofpacket    => id_router_031_src_endofpacket                                                 --          .endofpacket
		);

	id_router_032 : component NIOSIImicro_id_router_003
		port map (
			sink_ready         => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => pll_c0_clk,                                                                        --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                    -- clk_reset.reset
			src_ready          => id_router_032_src_ready,                                                           --       src.ready
			src_valid          => id_router_032_src_valid,                                                           --          .valid
			src_data           => id_router_032_src_data,                                                            --          .data
			src_channel        => id_router_032_src_channel,                                                         --          .channel
			src_startofpacket  => id_router_032_src_startofpacket,                                                   --          .startofpacket
			src_endofpacket    => id_router_032_src_endofpacket                                                      --          .endofpacket
		);

	limiter : component altera_merlin_traffic_limiter
		generic map (
			PKT_DEST_ID_H             => 93,
			PKT_DEST_ID_L             => 88,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			MAX_OUTSTANDING_RESPONSES => 9,
			PIPELINED                 => 0,
			ST_DATA_W                 => 104,
			ST_CHANNEL_W              => 33,
			VALID_WIDTH               => 33,
			ENFORCE_ORDER             => 1,
			PREVENT_HAZARDS           => 0,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32
		)
		port map (
			clk                    => pll_c0_clk,                     --       clk.clk
			reset                  => rst_controller_reset_out_reset, -- clk_reset.reset
			cmd_sink_ready         => addr_router_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_src_valid,          --          .valid
			cmd_sink_data          => addr_router_src_data,           --          .data
			cmd_sink_channel       => addr_router_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_cmd_src_ready,          --   cmd_src.ready
			cmd_src_data           => limiter_cmd_src_data,           --          .data
			cmd_src_channel        => limiter_cmd_src_channel,        --          .channel
			cmd_src_startofpacket  => limiter_cmd_src_startofpacket,  --          .startofpacket
			cmd_src_endofpacket    => limiter_cmd_src_endofpacket,    --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_rsp_src_ready,          --   rsp_src.ready
			rsp_src_valid          => limiter_rsp_src_valid,          --          .valid
			rsp_src_data           => limiter_rsp_src_data,           --          .data
			rsp_src_channel        => limiter_rsp_src_channel,        --          .channel
			rsp_src_startofpacket  => limiter_rsp_src_startofpacket,  --          .startofpacket
			rsp_src_endofpacket    => limiter_rsp_src_endofpacket,    --          .endofpacket
			cmd_src_valid          => limiter_cmd_valid_data          -- cmd_valid.data
		);

	burst_adapter : component altera_merlin_burst_adapter
		generic map (
			PKT_ADDR_H                => 42,
			PKT_ADDR_L                => 18,
			PKT_BEGIN_BURST           => 62,
			PKT_BYTE_CNT_H            => 51,
			PKT_BYTE_CNT_L            => 49,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_BURST_SIZE_H          => 57,
			PKT_BURST_SIZE_L          => 55,
			PKT_BURST_TYPE_H          => 59,
			PKT_BURST_TYPE_L          => 58,
			PKT_BURSTWRAP_H           => 54,
			PKT_BURSTWRAP_L           => 52,
			PKT_TRANS_COMPRESSED_READ => 43,
			PKT_TRANS_WRITE           => 45,
			PKT_TRANS_READ            => 46,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 86,
			ST_CHANNEL_W              => 33,
			OUT_BYTE_CNT_H            => 50,
			OUT_BURSTWRAP_H           => 54,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 3,
			BURSTWRAP_CONST_VALUE     => 3
		)
		port map (
			clk                   => pll_c0_clk,                          --       cr0.clk
			reset                 => rst_controller_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => width_adapter_src_valid,             --     sink0.valid
			sink0_data            => width_adapter_src_data,              --          .data
			sink0_channel         => width_adapter_src_channel,           --          .channel
			sink0_startofpacket   => width_adapter_src_startofpacket,     --          .startofpacket
			sink0_endofpacket     => width_adapter_src_endofpacket,       --          .endofpacket
			sink0_ready           => width_adapter_src_ready,             --          .ready
			source0_valid         => burst_adapter_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_source0_data,          --          .data
			source0_channel       => burst_adapter_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_source0_ready          --          .ready
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk        => pll_c0_clk,                     --       clk.clk
			reset_out  => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req  => open,                           -- (terminated)
			reset_in1  => '0',                            -- (terminated)
			reset_in2  => '0',                            -- (terminated)
			reset_in3  => '0',                            -- (terminated)
			reset_in4  => '0',                            -- (terminated)
			reset_in5  => '0',                            -- (terminated)
			reset_in6  => '0',                            -- (terminated)
			reset_in7  => '0',                            -- (terminated)
			reset_in8  => '0',                            -- (terminated)
			reset_in9  => '0',                            -- (terminated)
			reset_in10 => '0',                            -- (terminated)
			reset_in11 => '0',                            -- (terminated)
			reset_in12 => '0',                            -- (terminated)
			reset_in13 => '0',                            -- (terminated)
			reset_in14 => '0',                            -- (terminated)
			reset_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk        => clk_50_clk,                         --       clk.clk
			reset_out  => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req  => open,                               -- (terminated)
			reset_in1  => '0',                                -- (terminated)
			reset_in2  => '0',                                -- (terminated)
			reset_in3  => '0',                                -- (terminated)
			reset_in4  => '0',                                -- (terminated)
			reset_in5  => '0',                                -- (terminated)
			reset_in6  => '0',                                -- (terminated)
			reset_in7  => '0',                                -- (terminated)
			reset_in8  => '0',                                -- (terminated)
			reset_in9  => '0',                                -- (terminated)
			reset_in10 => '0',                                -- (terminated)
			reset_in11 => '0',                                -- (terminated)
			reset_in12 => '0',                                -- (terminated)
			reset_in13 => '0',                                -- (terminated)
			reset_in14 => '0',                                -- (terminated)
			reset_in15 => '0'                                 -- (terminated)
		);

	cmd_xbar_demux : component NIOSIImicro_cmd_xbar_demux
		port map (
			clk                => pll_c0_clk,                        --        clk.clk
			reset              => rst_controller_reset_out_reset,    --  clk_reset.reset
			sink_ready         => limiter_cmd_src_ready,             --       sink.ready
			sink_channel       => limiter_cmd_src_channel,           --           .channel
			sink_data          => limiter_cmd_src_data,              --           .data
			sink_startofpacket => limiter_cmd_src_startofpacket,     --           .startofpacket
			sink_endofpacket   => limiter_cmd_src_endofpacket,       --           .endofpacket
			sink_valid         => limiter_cmd_valid_data,            -- sink_valid.data
			src0_ready         => cmd_xbar_demux_src0_ready,         --       src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,         --           .valid
			src0_data          => cmd_xbar_demux_src0_data,          --           .data
			src0_channel       => cmd_xbar_demux_src0_channel,       --           .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket, --           .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,   --           .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,         --       src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,         --           .valid
			src1_data          => cmd_xbar_demux_src1_data,          --           .data
			src1_channel       => cmd_xbar_demux_src1_channel,       --           .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket, --           .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket,   --           .endofpacket
			src2_ready         => cmd_xbar_demux_src2_ready,         --       src2.ready
			src2_valid         => cmd_xbar_demux_src2_valid,         --           .valid
			src2_data          => cmd_xbar_demux_src2_data,          --           .data
			src2_channel       => cmd_xbar_demux_src2_channel,       --           .channel
			src2_startofpacket => cmd_xbar_demux_src2_startofpacket, --           .startofpacket
			src2_endofpacket   => cmd_xbar_demux_src2_endofpacket    --           .endofpacket
		);

	cmd_xbar_demux_001 : component NIOSIImicro_cmd_xbar_demux_001
		port map (
			clk                 => pll_c0_clk,                             --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			sink_ready          => addr_router_001_src_ready,              --      sink.ready
			sink_channel        => addr_router_001_src_channel,            --          .channel
			sink_data           => addr_router_001_src_data,               --          .data
			sink_startofpacket  => addr_router_001_src_startofpacket,      --          .startofpacket
			sink_endofpacket    => addr_router_001_src_endofpacket,        --          .endofpacket
			sink_valid(0)       => addr_router_001_src_valid,              --          .valid
			src0_ready          => cmd_xbar_demux_001_src0_ready,          --      src0.ready
			src0_valid          => cmd_xbar_demux_001_src0_valid,          --          .valid
			src0_data           => cmd_xbar_demux_001_src0_data,           --          .data
			src0_channel        => cmd_xbar_demux_001_src0_channel,        --          .channel
			src0_startofpacket  => cmd_xbar_demux_001_src0_startofpacket,  --          .startofpacket
			src0_endofpacket    => cmd_xbar_demux_001_src0_endofpacket,    --          .endofpacket
			src1_ready          => cmd_xbar_demux_001_src1_ready,          --      src1.ready
			src1_valid          => cmd_xbar_demux_001_src1_valid,          --          .valid
			src1_data           => cmd_xbar_demux_001_src1_data,           --          .data
			src1_channel        => cmd_xbar_demux_001_src1_channel,        --          .channel
			src1_startofpacket  => cmd_xbar_demux_001_src1_startofpacket,  --          .startofpacket
			src1_endofpacket    => cmd_xbar_demux_001_src1_endofpacket,    --          .endofpacket
			src2_ready          => cmd_xbar_demux_001_src2_ready,          --      src2.ready
			src2_valid          => cmd_xbar_demux_001_src2_valid,          --          .valid
			src2_data           => cmd_xbar_demux_001_src2_data,           --          .data
			src2_channel        => cmd_xbar_demux_001_src2_channel,        --          .channel
			src2_startofpacket  => cmd_xbar_demux_001_src2_startofpacket,  --          .startofpacket
			src2_endofpacket    => cmd_xbar_demux_001_src2_endofpacket,    --          .endofpacket
			src3_ready          => cmd_xbar_demux_001_src3_ready,          --      src3.ready
			src3_valid          => cmd_xbar_demux_001_src3_valid,          --          .valid
			src3_data           => cmd_xbar_demux_001_src3_data,           --          .data
			src3_channel        => cmd_xbar_demux_001_src3_channel,        --          .channel
			src3_startofpacket  => cmd_xbar_demux_001_src3_startofpacket,  --          .startofpacket
			src3_endofpacket    => cmd_xbar_demux_001_src3_endofpacket,    --          .endofpacket
			src4_ready          => cmd_xbar_demux_001_src4_ready,          --      src4.ready
			src4_valid          => cmd_xbar_demux_001_src4_valid,          --          .valid
			src4_data           => cmd_xbar_demux_001_src4_data,           --          .data
			src4_channel        => cmd_xbar_demux_001_src4_channel,        --          .channel
			src4_startofpacket  => cmd_xbar_demux_001_src4_startofpacket,  --          .startofpacket
			src4_endofpacket    => cmd_xbar_demux_001_src4_endofpacket,    --          .endofpacket
			src5_ready          => cmd_xbar_demux_001_src5_ready,          --      src5.ready
			src5_valid          => cmd_xbar_demux_001_src5_valid,          --          .valid
			src5_data           => cmd_xbar_demux_001_src5_data,           --          .data
			src5_channel        => cmd_xbar_demux_001_src5_channel,        --          .channel
			src5_startofpacket  => cmd_xbar_demux_001_src5_startofpacket,  --          .startofpacket
			src5_endofpacket    => cmd_xbar_demux_001_src5_endofpacket,    --          .endofpacket
			src6_ready          => cmd_xbar_demux_001_src6_ready,          --      src6.ready
			src6_valid          => cmd_xbar_demux_001_src6_valid,          --          .valid
			src6_data           => cmd_xbar_demux_001_src6_data,           --          .data
			src6_channel        => cmd_xbar_demux_001_src6_channel,        --          .channel
			src6_startofpacket  => cmd_xbar_demux_001_src6_startofpacket,  --          .startofpacket
			src6_endofpacket    => cmd_xbar_demux_001_src6_endofpacket,    --          .endofpacket
			src7_ready          => cmd_xbar_demux_001_src7_ready,          --      src7.ready
			src7_valid          => cmd_xbar_demux_001_src7_valid,          --          .valid
			src7_data           => cmd_xbar_demux_001_src7_data,           --          .data
			src7_channel        => cmd_xbar_demux_001_src7_channel,        --          .channel
			src7_startofpacket  => cmd_xbar_demux_001_src7_startofpacket,  --          .startofpacket
			src7_endofpacket    => cmd_xbar_demux_001_src7_endofpacket,    --          .endofpacket
			src8_ready          => cmd_xbar_demux_001_src8_ready,          --      src8.ready
			src8_valid          => cmd_xbar_demux_001_src8_valid,          --          .valid
			src8_data           => cmd_xbar_demux_001_src8_data,           --          .data
			src8_channel        => cmd_xbar_demux_001_src8_channel,        --          .channel
			src8_startofpacket  => cmd_xbar_demux_001_src8_startofpacket,  --          .startofpacket
			src8_endofpacket    => cmd_xbar_demux_001_src8_endofpacket,    --          .endofpacket
			src9_ready          => cmd_xbar_demux_001_src9_ready,          --      src9.ready
			src9_valid          => cmd_xbar_demux_001_src9_valid,          --          .valid
			src9_data           => cmd_xbar_demux_001_src9_data,           --          .data
			src9_channel        => cmd_xbar_demux_001_src9_channel,        --          .channel
			src9_startofpacket  => cmd_xbar_demux_001_src9_startofpacket,  --          .startofpacket
			src9_endofpacket    => cmd_xbar_demux_001_src9_endofpacket,    --          .endofpacket
			src10_ready         => cmd_xbar_demux_001_src10_ready,         --     src10.ready
			src10_valid         => cmd_xbar_demux_001_src10_valid,         --          .valid
			src10_data          => cmd_xbar_demux_001_src10_data,          --          .data
			src10_channel       => cmd_xbar_demux_001_src10_channel,       --          .channel
			src10_startofpacket => cmd_xbar_demux_001_src10_startofpacket, --          .startofpacket
			src10_endofpacket   => cmd_xbar_demux_001_src10_endofpacket,   --          .endofpacket
			src11_ready         => cmd_xbar_demux_001_src11_ready,         --     src11.ready
			src11_valid         => cmd_xbar_demux_001_src11_valid,         --          .valid
			src11_data          => cmd_xbar_demux_001_src11_data,          --          .data
			src11_channel       => cmd_xbar_demux_001_src11_channel,       --          .channel
			src11_startofpacket => cmd_xbar_demux_001_src11_startofpacket, --          .startofpacket
			src11_endofpacket   => cmd_xbar_demux_001_src11_endofpacket,   --          .endofpacket
			src12_ready         => cmd_xbar_demux_001_src12_ready,         --     src12.ready
			src12_valid         => cmd_xbar_demux_001_src12_valid,         --          .valid
			src12_data          => cmd_xbar_demux_001_src12_data,          --          .data
			src12_channel       => cmd_xbar_demux_001_src12_channel,       --          .channel
			src12_startofpacket => cmd_xbar_demux_001_src12_startofpacket, --          .startofpacket
			src12_endofpacket   => cmd_xbar_demux_001_src12_endofpacket,   --          .endofpacket
			src13_ready         => cmd_xbar_demux_001_src13_ready,         --     src13.ready
			src13_valid         => cmd_xbar_demux_001_src13_valid,         --          .valid
			src13_data          => cmd_xbar_demux_001_src13_data,          --          .data
			src13_channel       => cmd_xbar_demux_001_src13_channel,       --          .channel
			src13_startofpacket => cmd_xbar_demux_001_src13_startofpacket, --          .startofpacket
			src13_endofpacket   => cmd_xbar_demux_001_src13_endofpacket,   --          .endofpacket
			src14_ready         => cmd_xbar_demux_001_src14_ready,         --     src14.ready
			src14_valid         => cmd_xbar_demux_001_src14_valid,         --          .valid
			src14_data          => cmd_xbar_demux_001_src14_data,          --          .data
			src14_channel       => cmd_xbar_demux_001_src14_channel,       --          .channel
			src14_startofpacket => cmd_xbar_demux_001_src14_startofpacket, --          .startofpacket
			src14_endofpacket   => cmd_xbar_demux_001_src14_endofpacket,   --          .endofpacket
			src15_ready         => cmd_xbar_demux_001_src15_ready,         --     src15.ready
			src15_valid         => cmd_xbar_demux_001_src15_valid,         --          .valid
			src15_data          => cmd_xbar_demux_001_src15_data,          --          .data
			src15_channel       => cmd_xbar_demux_001_src15_channel,       --          .channel
			src15_startofpacket => cmd_xbar_demux_001_src15_startofpacket, --          .startofpacket
			src15_endofpacket   => cmd_xbar_demux_001_src15_endofpacket,   --          .endofpacket
			src16_ready         => cmd_xbar_demux_001_src16_ready,         --     src16.ready
			src16_valid         => cmd_xbar_demux_001_src16_valid,         --          .valid
			src16_data          => cmd_xbar_demux_001_src16_data,          --          .data
			src16_channel       => cmd_xbar_demux_001_src16_channel,       --          .channel
			src16_startofpacket => cmd_xbar_demux_001_src16_startofpacket, --          .startofpacket
			src16_endofpacket   => cmd_xbar_demux_001_src16_endofpacket,   --          .endofpacket
			src17_ready         => cmd_xbar_demux_001_src17_ready,         --     src17.ready
			src17_valid         => cmd_xbar_demux_001_src17_valid,         --          .valid
			src17_data          => cmd_xbar_demux_001_src17_data,          --          .data
			src17_channel       => cmd_xbar_demux_001_src17_channel,       --          .channel
			src17_startofpacket => cmd_xbar_demux_001_src17_startofpacket, --          .startofpacket
			src17_endofpacket   => cmd_xbar_demux_001_src17_endofpacket,   --          .endofpacket
			src18_ready         => cmd_xbar_demux_001_src18_ready,         --     src18.ready
			src18_valid         => cmd_xbar_demux_001_src18_valid,         --          .valid
			src18_data          => cmd_xbar_demux_001_src18_data,          --          .data
			src18_channel       => cmd_xbar_demux_001_src18_channel,       --          .channel
			src18_startofpacket => cmd_xbar_demux_001_src18_startofpacket, --          .startofpacket
			src18_endofpacket   => cmd_xbar_demux_001_src18_endofpacket,   --          .endofpacket
			src19_ready         => cmd_xbar_demux_001_src19_ready,         --     src19.ready
			src19_valid         => cmd_xbar_demux_001_src19_valid,         --          .valid
			src19_data          => cmd_xbar_demux_001_src19_data,          --          .data
			src19_channel       => cmd_xbar_demux_001_src19_channel,       --          .channel
			src19_startofpacket => cmd_xbar_demux_001_src19_startofpacket, --          .startofpacket
			src19_endofpacket   => cmd_xbar_demux_001_src19_endofpacket,   --          .endofpacket
			src20_ready         => cmd_xbar_demux_001_src20_ready,         --     src20.ready
			src20_valid         => cmd_xbar_demux_001_src20_valid,         --          .valid
			src20_data          => cmd_xbar_demux_001_src20_data,          --          .data
			src20_channel       => cmd_xbar_demux_001_src20_channel,       --          .channel
			src20_startofpacket => cmd_xbar_demux_001_src20_startofpacket, --          .startofpacket
			src20_endofpacket   => cmd_xbar_demux_001_src20_endofpacket,   --          .endofpacket
			src21_ready         => cmd_xbar_demux_001_src21_ready,         --     src21.ready
			src21_valid         => cmd_xbar_demux_001_src21_valid,         --          .valid
			src21_data          => cmd_xbar_demux_001_src21_data,          --          .data
			src21_channel       => cmd_xbar_demux_001_src21_channel,       --          .channel
			src21_startofpacket => cmd_xbar_demux_001_src21_startofpacket, --          .startofpacket
			src21_endofpacket   => cmd_xbar_demux_001_src21_endofpacket,   --          .endofpacket
			src22_ready         => cmd_xbar_demux_001_src22_ready,         --     src22.ready
			src22_valid         => cmd_xbar_demux_001_src22_valid,         --          .valid
			src22_data          => cmd_xbar_demux_001_src22_data,          --          .data
			src22_channel       => cmd_xbar_demux_001_src22_channel,       --          .channel
			src22_startofpacket => cmd_xbar_demux_001_src22_startofpacket, --          .startofpacket
			src22_endofpacket   => cmd_xbar_demux_001_src22_endofpacket,   --          .endofpacket
			src23_ready         => cmd_xbar_demux_001_src23_ready,         --     src23.ready
			src23_valid         => cmd_xbar_demux_001_src23_valid,         --          .valid
			src23_data          => cmd_xbar_demux_001_src23_data,          --          .data
			src23_channel       => cmd_xbar_demux_001_src23_channel,       --          .channel
			src23_startofpacket => cmd_xbar_demux_001_src23_startofpacket, --          .startofpacket
			src23_endofpacket   => cmd_xbar_demux_001_src23_endofpacket,   --          .endofpacket
			src24_ready         => cmd_xbar_demux_001_src24_ready,         --     src24.ready
			src24_valid         => cmd_xbar_demux_001_src24_valid,         --          .valid
			src24_data          => cmd_xbar_demux_001_src24_data,          --          .data
			src24_channel       => cmd_xbar_demux_001_src24_channel,       --          .channel
			src24_startofpacket => cmd_xbar_demux_001_src24_startofpacket, --          .startofpacket
			src24_endofpacket   => cmd_xbar_demux_001_src24_endofpacket,   --          .endofpacket
			src25_ready         => cmd_xbar_demux_001_src25_ready,         --     src25.ready
			src25_valid         => cmd_xbar_demux_001_src25_valid,         --          .valid
			src25_data          => cmd_xbar_demux_001_src25_data,          --          .data
			src25_channel       => cmd_xbar_demux_001_src25_channel,       --          .channel
			src25_startofpacket => cmd_xbar_demux_001_src25_startofpacket, --          .startofpacket
			src25_endofpacket   => cmd_xbar_demux_001_src25_endofpacket,   --          .endofpacket
			src26_ready         => cmd_xbar_demux_001_src26_ready,         --     src26.ready
			src26_valid         => cmd_xbar_demux_001_src26_valid,         --          .valid
			src26_data          => cmd_xbar_demux_001_src26_data,          --          .data
			src26_channel       => cmd_xbar_demux_001_src26_channel,       --          .channel
			src26_startofpacket => cmd_xbar_demux_001_src26_startofpacket, --          .startofpacket
			src26_endofpacket   => cmd_xbar_demux_001_src26_endofpacket,   --          .endofpacket
			src27_ready         => cmd_xbar_demux_001_src27_ready,         --     src27.ready
			src27_valid         => cmd_xbar_demux_001_src27_valid,         --          .valid
			src27_data          => cmd_xbar_demux_001_src27_data,          --          .data
			src27_channel       => cmd_xbar_demux_001_src27_channel,       --          .channel
			src27_startofpacket => cmd_xbar_demux_001_src27_startofpacket, --          .startofpacket
			src27_endofpacket   => cmd_xbar_demux_001_src27_endofpacket,   --          .endofpacket
			src28_ready         => cmd_xbar_demux_001_src28_ready,         --     src28.ready
			src28_valid         => cmd_xbar_demux_001_src28_valid,         --          .valid
			src28_data          => cmd_xbar_demux_001_src28_data,          --          .data
			src28_channel       => cmd_xbar_demux_001_src28_channel,       --          .channel
			src28_startofpacket => cmd_xbar_demux_001_src28_startofpacket, --          .startofpacket
			src28_endofpacket   => cmd_xbar_demux_001_src28_endofpacket,   --          .endofpacket
			src29_ready         => cmd_xbar_demux_001_src29_ready,         --     src29.ready
			src29_valid         => cmd_xbar_demux_001_src29_valid,         --          .valid
			src29_data          => cmd_xbar_demux_001_src29_data,          --          .data
			src29_channel       => cmd_xbar_demux_001_src29_channel,       --          .channel
			src29_startofpacket => cmd_xbar_demux_001_src29_startofpacket, --          .startofpacket
			src29_endofpacket   => cmd_xbar_demux_001_src29_endofpacket,   --          .endofpacket
			src30_ready         => cmd_xbar_demux_001_src30_ready,         --     src30.ready
			src30_valid         => cmd_xbar_demux_001_src30_valid,         --          .valid
			src30_data          => cmd_xbar_demux_001_src30_data,          --          .data
			src30_channel       => cmd_xbar_demux_001_src30_channel,       --          .channel
			src30_startofpacket => cmd_xbar_demux_001_src30_startofpacket, --          .startofpacket
			src30_endofpacket   => cmd_xbar_demux_001_src30_endofpacket,   --          .endofpacket
			src31_ready         => cmd_xbar_demux_001_src31_ready,         --     src31.ready
			src31_valid         => cmd_xbar_demux_001_src31_valid,         --          .valid
			src31_data          => cmd_xbar_demux_001_src31_data,          --          .data
			src31_channel       => cmd_xbar_demux_001_src31_channel,       --          .channel
			src31_startofpacket => cmd_xbar_demux_001_src31_startofpacket, --          .startofpacket
			src31_endofpacket   => cmd_xbar_demux_001_src31_endofpacket,   --          .endofpacket
			src32_ready         => cmd_xbar_demux_001_src32_ready,         --     src32.ready
			src32_valid         => cmd_xbar_demux_001_src32_valid,         --          .valid
			src32_data          => cmd_xbar_demux_001_src32_data,          --          .data
			src32_channel       => cmd_xbar_demux_001_src32_channel,       --          .channel
			src32_startofpacket => cmd_xbar_demux_001_src32_startofpacket, --          .startofpacket
			src32_endofpacket   => cmd_xbar_demux_001_src32_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux : component NIOSIImicro_cmd_xbar_mux
		port map (
			clk                 => pll_c0_clk,                            --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component NIOSIImicro_cmd_xbar_mux
		port map (
			clk                 => pll_c0_clk,                            --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_002 : component NIOSIImicro_cmd_xbar_mux
		port map (
			clk                 => pll_c0_clk,                            --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_002_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_002_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_002_src_data,             --          .data
			src_channel         => cmd_xbar_mux_002_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_002_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_002_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src2_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src2_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src2_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src2_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src2_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src2_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src2_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src2_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src2_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src2_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src2_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux : component NIOSIImicro_rsp_xbar_demux
		port map (
			clk                => pll_c0_clk,                        --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_src_ready,               --      sink.ready
			sink_channel       => id_router_src_channel,             --          .channel
			sink_data          => id_router_src_data,                --          .data
			sink_startofpacket => id_router_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_001 : component NIOSIImicro_rsp_xbar_demux
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => width_adapter_001_src_ready,           --      sink.ready
			sink_channel       => width_adapter_001_src_channel,         --          .channel
			sink_data          => width_adapter_001_src_data,            --          .data
			sink_startofpacket => width_adapter_001_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_001_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_001_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component NIOSIImicro_rsp_xbar_demux
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_002_src_ready,               --      sink.ready
			sink_channel       => id_router_002_src_channel,             --          .channel
			sink_data          => id_router_002_src_data,                --          .data
			sink_startofpacket => id_router_002_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_002_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_002_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_002_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_002_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_002_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_002_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_002_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => clk_50_clk,                            --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_003_src_ready,               --      sink.ready
			sink_channel       => id_router_003_src_channel,             --          .channel
			sink_data          => id_router_003_src_data,                --          .data
			sink_startofpacket => id_router_003_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_003_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_003_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,               --      sink.ready
			sink_channel       => id_router_004_src_channel,             --          .channel
			sink_data          => id_router_004_src_data,                --          .data
			sink_startofpacket => id_router_004_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,               --      sink.ready
			sink_channel       => id_router_005_src_channel,             --          .channel
			sink_data          => id_router_005_src_data,                --          .data
			sink_startofpacket => id_router_005_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,               --      sink.ready
			sink_channel       => id_router_006_src_channel,             --          .channel
			sink_data          => id_router_006_src_data,                --          .data
			sink_startofpacket => id_router_006_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_007 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_007_src_ready,               --      sink.ready
			sink_channel       => id_router_007_src_channel,             --          .channel
			sink_data          => id_router_007_src_data,                --          .data
			sink_startofpacket => id_router_007_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_007_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_007_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_008 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_008_src_ready,               --      sink.ready
			sink_channel       => id_router_008_src_channel,             --          .channel
			sink_data          => id_router_008_src_data,                --          .data
			sink_startofpacket => id_router_008_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_008_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_008_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_008_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_008_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_008_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_009 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_009_src_ready,               --      sink.ready
			sink_channel       => id_router_009_src_channel,             --          .channel
			sink_data          => id_router_009_src_data,                --          .data
			sink_startofpacket => id_router_009_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_009_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_009_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_009_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_009_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_009_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_010 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_010_src_ready,               --      sink.ready
			sink_channel       => id_router_010_src_channel,             --          .channel
			sink_data          => id_router_010_src_data,                --          .data
			sink_startofpacket => id_router_010_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_010_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_010_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_010_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_010_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_010_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_011 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_011_src_ready,               --      sink.ready
			sink_channel       => id_router_011_src_channel,             --          .channel
			sink_data          => id_router_011_src_data,                --          .data
			sink_startofpacket => id_router_011_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_011_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_011_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_011_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_011_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_011_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_012 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_012_src_ready,               --      sink.ready
			sink_channel       => id_router_012_src_channel,             --          .channel
			sink_data          => id_router_012_src_data,                --          .data
			sink_startofpacket => id_router_012_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_012_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_012_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_012_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_012_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_012_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_013 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_013_src_ready,               --      sink.ready
			sink_channel       => id_router_013_src_channel,             --          .channel
			sink_data          => id_router_013_src_data,                --          .data
			sink_startofpacket => id_router_013_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_013_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_013_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_013_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_013_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_013_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_014 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_014_src_ready,               --      sink.ready
			sink_channel       => id_router_014_src_channel,             --          .channel
			sink_data          => id_router_014_src_data,                --          .data
			sink_startofpacket => id_router_014_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_014_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_014_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_014_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_014_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_014_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_014_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_014_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_014_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_015 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_015_src_ready,               --      sink.ready
			sink_channel       => id_router_015_src_channel,             --          .channel
			sink_data          => id_router_015_src_data,                --          .data
			sink_startofpacket => id_router_015_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_015_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_015_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_015_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_015_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_015_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_015_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_015_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_015_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_016 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_016_src_ready,               --      sink.ready
			sink_channel       => id_router_016_src_channel,             --          .channel
			sink_data          => id_router_016_src_data,                --          .data
			sink_startofpacket => id_router_016_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_016_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_016_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_016_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_016_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_016_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_016_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_016_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_016_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_017 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_017_src_ready,               --      sink.ready
			sink_channel       => id_router_017_src_channel,             --          .channel
			sink_data          => id_router_017_src_data,                --          .data
			sink_startofpacket => id_router_017_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_017_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_017_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_017_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_017_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_017_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_017_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_017_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_017_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_018 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_018_src_ready,               --      sink.ready
			sink_channel       => id_router_018_src_channel,             --          .channel
			sink_data          => id_router_018_src_data,                --          .data
			sink_startofpacket => id_router_018_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_018_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_018_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_018_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_018_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_018_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_018_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_018_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_018_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_019 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_019_src_ready,               --      sink.ready
			sink_channel       => id_router_019_src_channel,             --          .channel
			sink_data          => id_router_019_src_data,                --          .data
			sink_startofpacket => id_router_019_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_019_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_019_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_019_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_019_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_019_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_019_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_019_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_019_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_020 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_020_src_ready,               --      sink.ready
			sink_channel       => id_router_020_src_channel,             --          .channel
			sink_data          => id_router_020_src_data,                --          .data
			sink_startofpacket => id_router_020_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_020_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_020_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_020_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_020_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_020_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_020_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_020_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_020_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_021 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_021_src_ready,               --      sink.ready
			sink_channel       => id_router_021_src_channel,             --          .channel
			sink_data          => id_router_021_src_data,                --          .data
			sink_startofpacket => id_router_021_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_021_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_021_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_021_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_021_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_021_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_021_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_021_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_021_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_022 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_022_src_ready,               --      sink.ready
			sink_channel       => id_router_022_src_channel,             --          .channel
			sink_data          => id_router_022_src_data,                --          .data
			sink_startofpacket => id_router_022_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_022_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_022_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_022_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_022_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_022_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_022_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_022_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_022_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_023 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_023_src_ready,               --      sink.ready
			sink_channel       => id_router_023_src_channel,             --          .channel
			sink_data          => id_router_023_src_data,                --          .data
			sink_startofpacket => id_router_023_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_023_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_023_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_023_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_023_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_023_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_023_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_023_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_023_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_024 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_024_src_ready,               --      sink.ready
			sink_channel       => id_router_024_src_channel,             --          .channel
			sink_data          => id_router_024_src_data,                --          .data
			sink_startofpacket => id_router_024_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_024_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_024_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_024_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_024_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_024_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_024_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_024_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_024_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_025 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_025_src_ready,               --      sink.ready
			sink_channel       => id_router_025_src_channel,             --          .channel
			sink_data          => id_router_025_src_data,                --          .data
			sink_startofpacket => id_router_025_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_025_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_025_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_025_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_025_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_025_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_025_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_025_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_025_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_026 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_026_src_ready,               --      sink.ready
			sink_channel       => id_router_026_src_channel,             --          .channel
			sink_data          => id_router_026_src_data,                --          .data
			sink_startofpacket => id_router_026_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_026_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_026_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_026_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_026_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_026_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_026_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_026_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_026_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_027 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_027_src_ready,               --      sink.ready
			sink_channel       => id_router_027_src_channel,             --          .channel
			sink_data          => id_router_027_src_data,                --          .data
			sink_startofpacket => id_router_027_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_027_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_027_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_027_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_027_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_027_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_027_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_027_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_027_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_028 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_028_src_ready,               --      sink.ready
			sink_channel       => id_router_028_src_channel,             --          .channel
			sink_data          => id_router_028_src_data,                --          .data
			sink_startofpacket => id_router_028_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_028_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_028_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_028_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_028_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_028_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_028_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_028_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_028_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_029 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_029_src_ready,               --      sink.ready
			sink_channel       => id_router_029_src_channel,             --          .channel
			sink_data          => id_router_029_src_data,                --          .data
			sink_startofpacket => id_router_029_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_029_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_029_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_029_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_029_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_029_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_029_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_029_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_029_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_030 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_030_src_ready,               --      sink.ready
			sink_channel       => id_router_030_src_channel,             --          .channel
			sink_data          => id_router_030_src_data,                --          .data
			sink_startofpacket => id_router_030_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_030_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_030_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_030_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_030_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_030_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_030_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_030_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_030_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_031 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_031_src_ready,               --      sink.ready
			sink_channel       => id_router_031_src_channel,             --          .channel
			sink_data          => id_router_031_src_data,                --          .data
			sink_startofpacket => id_router_031_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_031_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_031_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_031_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_031_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_031_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_031_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_031_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_031_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_032 : component NIOSIImicro_rsp_xbar_demux_003
		port map (
			clk                => pll_c0_clk,                            --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_032_src_ready,               --      sink.ready
			sink_channel       => id_router_032_src_channel,             --          .channel
			sink_data          => id_router_032_src_data,                --          .data
			sink_startofpacket => id_router_032_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_032_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_032_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_032_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_032_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_032_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_032_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_032_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_032_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component NIOSIImicro_rsp_xbar_mux
		port map (
			clk                 => pll_c0_clk,                            --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,                --          .valid
			src_data            => rsp_xbar_mux_src_data,                 --          .data
			src_channel         => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_002_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_001 : component NIOSIImicro_rsp_xbar_mux_001
		port map (
			clk                  => pll_c0_clk,                            --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready            => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid            => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data             => rsp_xbar_mux_001_src_data,             --          .data
			src_channel          => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket    => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket      => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready          => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid          => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel        => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data           => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket  => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket    => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready          => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid          => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel        => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data           => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket  => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket    => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			sink2_ready          => rsp_xbar_demux_002_src1_ready,         --     sink2.ready
			sink2_valid          => rsp_xbar_demux_002_src1_valid,         --          .valid
			sink2_channel        => rsp_xbar_demux_002_src1_channel,       --          .channel
			sink2_data           => rsp_xbar_demux_002_src1_data,          --          .data
			sink2_startofpacket  => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			sink2_endofpacket    => rsp_xbar_demux_002_src1_endofpacket,   --          .endofpacket
			sink3_ready          => crosser_001_out_ready,                 --     sink3.ready
			sink3_valid          => crosser_001_out_valid,                 --          .valid
			sink3_channel        => crosser_001_out_channel,               --          .channel
			sink3_data           => crosser_001_out_data,                  --          .data
			sink3_startofpacket  => crosser_001_out_startofpacket,         --          .startofpacket
			sink3_endofpacket    => crosser_001_out_endofpacket,           --          .endofpacket
			sink4_ready          => rsp_xbar_demux_004_src0_ready,         --     sink4.ready
			sink4_valid          => rsp_xbar_demux_004_src0_valid,         --          .valid
			sink4_channel        => rsp_xbar_demux_004_src0_channel,       --          .channel
			sink4_data           => rsp_xbar_demux_004_src0_data,          --          .data
			sink4_startofpacket  => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink4_endofpacket    => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			sink5_ready          => rsp_xbar_demux_005_src0_ready,         --     sink5.ready
			sink5_valid          => rsp_xbar_demux_005_src0_valid,         --          .valid
			sink5_channel        => rsp_xbar_demux_005_src0_channel,       --          .channel
			sink5_data           => rsp_xbar_demux_005_src0_data,          --          .data
			sink5_startofpacket  => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			sink5_endofpacket    => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			sink6_ready          => rsp_xbar_demux_006_src0_ready,         --     sink6.ready
			sink6_valid          => rsp_xbar_demux_006_src0_valid,         --          .valid
			sink6_channel        => rsp_xbar_demux_006_src0_channel,       --          .channel
			sink6_data           => rsp_xbar_demux_006_src0_data,          --          .data
			sink6_startofpacket  => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink6_endofpacket    => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			sink7_ready          => rsp_xbar_demux_007_src0_ready,         --     sink7.ready
			sink7_valid          => rsp_xbar_demux_007_src0_valid,         --          .valid
			sink7_channel        => rsp_xbar_demux_007_src0_channel,       --          .channel
			sink7_data           => rsp_xbar_demux_007_src0_data,          --          .data
			sink7_startofpacket  => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			sink7_endofpacket    => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			sink8_ready          => rsp_xbar_demux_008_src0_ready,         --     sink8.ready
			sink8_valid          => rsp_xbar_demux_008_src0_valid,         --          .valid
			sink8_channel        => rsp_xbar_demux_008_src0_channel,       --          .channel
			sink8_data           => rsp_xbar_demux_008_src0_data,          --          .data
			sink8_startofpacket  => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			sink8_endofpacket    => rsp_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			sink9_ready          => rsp_xbar_demux_009_src0_ready,         --     sink9.ready
			sink9_valid          => rsp_xbar_demux_009_src0_valid,         --          .valid
			sink9_channel        => rsp_xbar_demux_009_src0_channel,       --          .channel
			sink9_data           => rsp_xbar_demux_009_src0_data,          --          .data
			sink9_startofpacket  => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			sink9_endofpacket    => rsp_xbar_demux_009_src0_endofpacket,   --          .endofpacket
			sink10_ready         => rsp_xbar_demux_010_src0_ready,         --    sink10.ready
			sink10_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			sink10_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			sink10_data          => rsp_xbar_demux_010_src0_data,          --          .data
			sink10_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			sink10_endofpacket   => rsp_xbar_demux_010_src0_endofpacket,   --          .endofpacket
			sink11_ready         => rsp_xbar_demux_011_src0_ready,         --    sink11.ready
			sink11_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			sink11_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			sink11_data          => rsp_xbar_demux_011_src0_data,          --          .data
			sink11_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			sink11_endofpacket   => rsp_xbar_demux_011_src0_endofpacket,   --          .endofpacket
			sink12_ready         => rsp_xbar_demux_012_src0_ready,         --    sink12.ready
			sink12_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			sink12_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			sink12_data          => rsp_xbar_demux_012_src0_data,          --          .data
			sink12_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			sink12_endofpacket   => rsp_xbar_demux_012_src0_endofpacket,   --          .endofpacket
			sink13_ready         => rsp_xbar_demux_013_src0_ready,         --    sink13.ready
			sink13_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			sink13_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			sink13_data          => rsp_xbar_demux_013_src0_data,          --          .data
			sink13_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			sink13_endofpacket   => rsp_xbar_demux_013_src0_endofpacket,   --          .endofpacket
			sink14_ready         => rsp_xbar_demux_014_src0_ready,         --    sink14.ready
			sink14_valid         => rsp_xbar_demux_014_src0_valid,         --          .valid
			sink14_channel       => rsp_xbar_demux_014_src0_channel,       --          .channel
			sink14_data          => rsp_xbar_demux_014_src0_data,          --          .data
			sink14_startofpacket => rsp_xbar_demux_014_src0_startofpacket, --          .startofpacket
			sink14_endofpacket   => rsp_xbar_demux_014_src0_endofpacket,   --          .endofpacket
			sink15_ready         => rsp_xbar_demux_015_src0_ready,         --    sink15.ready
			sink15_valid         => rsp_xbar_demux_015_src0_valid,         --          .valid
			sink15_channel       => rsp_xbar_demux_015_src0_channel,       --          .channel
			sink15_data          => rsp_xbar_demux_015_src0_data,          --          .data
			sink15_startofpacket => rsp_xbar_demux_015_src0_startofpacket, --          .startofpacket
			sink15_endofpacket   => rsp_xbar_demux_015_src0_endofpacket,   --          .endofpacket
			sink16_ready         => rsp_xbar_demux_016_src0_ready,         --    sink16.ready
			sink16_valid         => rsp_xbar_demux_016_src0_valid,         --          .valid
			sink16_channel       => rsp_xbar_demux_016_src0_channel,       --          .channel
			sink16_data          => rsp_xbar_demux_016_src0_data,          --          .data
			sink16_startofpacket => rsp_xbar_demux_016_src0_startofpacket, --          .startofpacket
			sink16_endofpacket   => rsp_xbar_demux_016_src0_endofpacket,   --          .endofpacket
			sink17_ready         => rsp_xbar_demux_017_src0_ready,         --    sink17.ready
			sink17_valid         => rsp_xbar_demux_017_src0_valid,         --          .valid
			sink17_channel       => rsp_xbar_demux_017_src0_channel,       --          .channel
			sink17_data          => rsp_xbar_demux_017_src0_data,          --          .data
			sink17_startofpacket => rsp_xbar_demux_017_src0_startofpacket, --          .startofpacket
			sink17_endofpacket   => rsp_xbar_demux_017_src0_endofpacket,   --          .endofpacket
			sink18_ready         => rsp_xbar_demux_018_src0_ready,         --    sink18.ready
			sink18_valid         => rsp_xbar_demux_018_src0_valid,         --          .valid
			sink18_channel       => rsp_xbar_demux_018_src0_channel,       --          .channel
			sink18_data          => rsp_xbar_demux_018_src0_data,          --          .data
			sink18_startofpacket => rsp_xbar_demux_018_src0_startofpacket, --          .startofpacket
			sink18_endofpacket   => rsp_xbar_demux_018_src0_endofpacket,   --          .endofpacket
			sink19_ready         => rsp_xbar_demux_019_src0_ready,         --    sink19.ready
			sink19_valid         => rsp_xbar_demux_019_src0_valid,         --          .valid
			sink19_channel       => rsp_xbar_demux_019_src0_channel,       --          .channel
			sink19_data          => rsp_xbar_demux_019_src0_data,          --          .data
			sink19_startofpacket => rsp_xbar_demux_019_src0_startofpacket, --          .startofpacket
			sink19_endofpacket   => rsp_xbar_demux_019_src0_endofpacket,   --          .endofpacket
			sink20_ready         => rsp_xbar_demux_020_src0_ready,         --    sink20.ready
			sink20_valid         => rsp_xbar_demux_020_src0_valid,         --          .valid
			sink20_channel       => rsp_xbar_demux_020_src0_channel,       --          .channel
			sink20_data          => rsp_xbar_demux_020_src0_data,          --          .data
			sink20_startofpacket => rsp_xbar_demux_020_src0_startofpacket, --          .startofpacket
			sink20_endofpacket   => rsp_xbar_demux_020_src0_endofpacket,   --          .endofpacket
			sink21_ready         => rsp_xbar_demux_021_src0_ready,         --    sink21.ready
			sink21_valid         => rsp_xbar_demux_021_src0_valid,         --          .valid
			sink21_channel       => rsp_xbar_demux_021_src0_channel,       --          .channel
			sink21_data          => rsp_xbar_demux_021_src0_data,          --          .data
			sink21_startofpacket => rsp_xbar_demux_021_src0_startofpacket, --          .startofpacket
			sink21_endofpacket   => rsp_xbar_demux_021_src0_endofpacket,   --          .endofpacket
			sink22_ready         => rsp_xbar_demux_022_src0_ready,         --    sink22.ready
			sink22_valid         => rsp_xbar_demux_022_src0_valid,         --          .valid
			sink22_channel       => rsp_xbar_demux_022_src0_channel,       --          .channel
			sink22_data          => rsp_xbar_demux_022_src0_data,          --          .data
			sink22_startofpacket => rsp_xbar_demux_022_src0_startofpacket, --          .startofpacket
			sink22_endofpacket   => rsp_xbar_demux_022_src0_endofpacket,   --          .endofpacket
			sink23_ready         => rsp_xbar_demux_023_src0_ready,         --    sink23.ready
			sink23_valid         => rsp_xbar_demux_023_src0_valid,         --          .valid
			sink23_channel       => rsp_xbar_demux_023_src0_channel,       --          .channel
			sink23_data          => rsp_xbar_demux_023_src0_data,          --          .data
			sink23_startofpacket => rsp_xbar_demux_023_src0_startofpacket, --          .startofpacket
			sink23_endofpacket   => rsp_xbar_demux_023_src0_endofpacket,   --          .endofpacket
			sink24_ready         => rsp_xbar_demux_024_src0_ready,         --    sink24.ready
			sink24_valid         => rsp_xbar_demux_024_src0_valid,         --          .valid
			sink24_channel       => rsp_xbar_demux_024_src0_channel,       --          .channel
			sink24_data          => rsp_xbar_demux_024_src0_data,          --          .data
			sink24_startofpacket => rsp_xbar_demux_024_src0_startofpacket, --          .startofpacket
			sink24_endofpacket   => rsp_xbar_demux_024_src0_endofpacket,   --          .endofpacket
			sink25_ready         => rsp_xbar_demux_025_src0_ready,         --    sink25.ready
			sink25_valid         => rsp_xbar_demux_025_src0_valid,         --          .valid
			sink25_channel       => rsp_xbar_demux_025_src0_channel,       --          .channel
			sink25_data          => rsp_xbar_demux_025_src0_data,          --          .data
			sink25_startofpacket => rsp_xbar_demux_025_src0_startofpacket, --          .startofpacket
			sink25_endofpacket   => rsp_xbar_demux_025_src0_endofpacket,   --          .endofpacket
			sink26_ready         => rsp_xbar_demux_026_src0_ready,         --    sink26.ready
			sink26_valid         => rsp_xbar_demux_026_src0_valid,         --          .valid
			sink26_channel       => rsp_xbar_demux_026_src0_channel,       --          .channel
			sink26_data          => rsp_xbar_demux_026_src0_data,          --          .data
			sink26_startofpacket => rsp_xbar_demux_026_src0_startofpacket, --          .startofpacket
			sink26_endofpacket   => rsp_xbar_demux_026_src0_endofpacket,   --          .endofpacket
			sink27_ready         => rsp_xbar_demux_027_src0_ready,         --    sink27.ready
			sink27_valid         => rsp_xbar_demux_027_src0_valid,         --          .valid
			sink27_channel       => rsp_xbar_demux_027_src0_channel,       --          .channel
			sink27_data          => rsp_xbar_demux_027_src0_data,          --          .data
			sink27_startofpacket => rsp_xbar_demux_027_src0_startofpacket, --          .startofpacket
			sink27_endofpacket   => rsp_xbar_demux_027_src0_endofpacket,   --          .endofpacket
			sink28_ready         => rsp_xbar_demux_028_src0_ready,         --    sink28.ready
			sink28_valid         => rsp_xbar_demux_028_src0_valid,         --          .valid
			sink28_channel       => rsp_xbar_demux_028_src0_channel,       --          .channel
			sink28_data          => rsp_xbar_demux_028_src0_data,          --          .data
			sink28_startofpacket => rsp_xbar_demux_028_src0_startofpacket, --          .startofpacket
			sink28_endofpacket   => rsp_xbar_demux_028_src0_endofpacket,   --          .endofpacket
			sink29_ready         => rsp_xbar_demux_029_src0_ready,         --    sink29.ready
			sink29_valid         => rsp_xbar_demux_029_src0_valid,         --          .valid
			sink29_channel       => rsp_xbar_demux_029_src0_channel,       --          .channel
			sink29_data          => rsp_xbar_demux_029_src0_data,          --          .data
			sink29_startofpacket => rsp_xbar_demux_029_src0_startofpacket, --          .startofpacket
			sink29_endofpacket   => rsp_xbar_demux_029_src0_endofpacket,   --          .endofpacket
			sink30_ready         => rsp_xbar_demux_030_src0_ready,         --    sink30.ready
			sink30_valid         => rsp_xbar_demux_030_src0_valid,         --          .valid
			sink30_channel       => rsp_xbar_demux_030_src0_channel,       --          .channel
			sink30_data          => rsp_xbar_demux_030_src0_data,          --          .data
			sink30_startofpacket => rsp_xbar_demux_030_src0_startofpacket, --          .startofpacket
			sink30_endofpacket   => rsp_xbar_demux_030_src0_endofpacket,   --          .endofpacket
			sink31_ready         => rsp_xbar_demux_031_src0_ready,         --    sink31.ready
			sink31_valid         => rsp_xbar_demux_031_src0_valid,         --          .valid
			sink31_channel       => rsp_xbar_demux_031_src0_channel,       --          .channel
			sink31_data          => rsp_xbar_demux_031_src0_data,          --          .data
			sink31_startofpacket => rsp_xbar_demux_031_src0_startofpacket, --          .startofpacket
			sink31_endofpacket   => rsp_xbar_demux_031_src0_endofpacket,   --          .endofpacket
			sink32_ready         => rsp_xbar_demux_032_src0_ready,         --    sink32.ready
			sink32_valid         => rsp_xbar_demux_032_src0_valid,         --          .valid
			sink32_channel       => rsp_xbar_demux_032_src0_channel,       --          .channel
			sink32_data          => rsp_xbar_demux_032_src0_data,          --          .data
			sink32_startofpacket => rsp_xbar_demux_032_src0_startofpacket, --          .startofpacket
			sink32_endofpacket   => rsp_xbar_demux_032_src0_endofpacket    --          .endofpacket
		);

	width_adapter : component niosiimicro_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 60,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 69,
			IN_PKT_BYTE_CNT_L             => 67,
			IN_PKT_TRANS_COMPRESSED_READ  => 61,
			IN_PKT_BURSTWRAP_H            => 72,
			IN_PKT_BURSTWRAP_L            => 70,
			IN_PKT_BURST_SIZE_H           => 75,
			IN_PKT_BURST_SIZE_L           => 73,
			IN_PKT_RESPONSE_STATUS_H      => 103,
			IN_PKT_RESPONSE_STATUS_L      => 102,
			IN_PKT_TRANS_EXCLUSIVE        => 66,
			IN_PKT_BURST_TYPE_H           => 77,
			IN_PKT_BURST_TYPE_L           => 76,
			IN_ST_DATA_W                  => 104,
			OUT_PKT_ADDR_H                => 42,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 51,
			OUT_PKT_BYTE_CNT_L            => 49,
			OUT_PKT_TRANS_COMPRESSED_READ => 43,
			OUT_PKT_BURST_SIZE_H          => 57,
			OUT_PKT_BURST_SIZE_L          => 55,
			OUT_PKT_RESPONSE_STATUS_H     => 85,
			OUT_PKT_RESPONSE_STATUS_L     => 84,
			OUT_PKT_TRANS_EXCLUSIVE       => 48,
			OUT_PKT_BURST_TYPE_H          => 59,
			OUT_PKT_BURST_TYPE_L          => 58,
			OUT_ST_DATA_W                 => 86,
			ST_CHANNEL_W                  => 33,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => pll_c0_clk,                         --       clk.clk
			reset                => rst_controller_reset_out_reset,     -- clk_reset.reset
			in_valid             => cmd_xbar_mux_001_src_valid,         --      sink.valid
			in_channel           => cmd_xbar_mux_001_src_channel,       --          .channel
			in_startofpacket     => cmd_xbar_mux_001_src_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_mux_001_src_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_mux_001_src_ready,         --          .ready
			in_data              => cmd_xbar_mux_001_src_data,          --          .data
			out_endofpacket      => width_adapter_src_endofpacket,      --       src.endofpacket
			out_data             => width_adapter_src_data,             --          .data
			out_channel          => width_adapter_src_channel,          --          .channel
			out_valid            => width_adapter_src_valid,            --          .valid
			out_ready            => width_adapter_src_ready,            --          .ready
			out_startofpacket    => width_adapter_src_startofpacket,    --          .startofpacket
			in_command_size_data => "000"                               -- (terminated)
		);

	width_adapter_001 : component niosiimicro_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 42,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 51,
			IN_PKT_BYTE_CNT_L             => 49,
			IN_PKT_TRANS_COMPRESSED_READ  => 43,
			IN_PKT_BURSTWRAP_H            => 54,
			IN_PKT_BURSTWRAP_L            => 52,
			IN_PKT_BURST_SIZE_H           => 57,
			IN_PKT_BURST_SIZE_L           => 55,
			IN_PKT_RESPONSE_STATUS_H      => 85,
			IN_PKT_RESPONSE_STATUS_L      => 84,
			IN_PKT_TRANS_EXCLUSIVE        => 48,
			IN_PKT_BURST_TYPE_H           => 59,
			IN_PKT_BURST_TYPE_L           => 58,
			IN_ST_DATA_W                  => 86,
			OUT_PKT_ADDR_H                => 60,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 69,
			OUT_PKT_BYTE_CNT_L            => 67,
			OUT_PKT_TRANS_COMPRESSED_READ => 61,
			OUT_PKT_BURST_SIZE_H          => 75,
			OUT_PKT_BURST_SIZE_L          => 73,
			OUT_PKT_RESPONSE_STATUS_H     => 103,
			OUT_PKT_RESPONSE_STATUS_L     => 102,
			OUT_PKT_TRANS_EXCLUSIVE       => 66,
			OUT_PKT_BURST_TYPE_H          => 77,
			OUT_PKT_BURST_TYPE_L          => 76,
			OUT_ST_DATA_W                 => 104,
			ST_CHANNEL_W                  => 33,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => pll_c0_clk,                          --       clk.clk
			reset                => rst_controller_reset_out_reset,      -- clk_reset.reset
			in_valid             => id_router_001_src_valid,             --      sink.valid
			in_channel           => id_router_001_src_channel,           --          .channel
			in_startofpacket     => id_router_001_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_001_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_001_src_ready,             --          .ready
			in_data              => id_router_001_src_data,              --          .data
			out_endofpacket      => width_adapter_001_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_001_src_data,          --          .data
			out_channel          => width_adapter_001_src_channel,       --          .channel
			out_valid            => width_adapter_001_src_valid,         --          .valid
			out_ready            => width_adapter_001_src_ready,         --          .ready
			out_startofpacket    => width_adapter_001_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	crosser : component altera_avalon_st_handshake_clock_crosser
		generic map (
			DATA_WIDTH          => 104,
			BITS_PER_SYMBOL     => 104,
			USE_PACKETS         => 1,
			USE_CHANNEL         => 1,
			CHANNEL_WIDTH       => 33,
			USE_ERROR           => 0,
			ERROR_WIDTH         => 1,
			VALID_SYNC_DEPTH    => 2,
			READY_SYNC_DEPTH    => 2,
			USE_OUTPUT_PIPELINE => 0
		)
		port map (
			in_clk            => pll_c0_clk,                            --        in_clk.clk
			in_reset          => rst_controller_reset_out_reset,        --  in_clk_reset.reset
			out_clk           => clk_50_clk,                            --       out_clk.clk
			out_reset         => rst_controller_001_reset_out_reset,    -- out_clk_reset.reset
			in_ready          => cmd_xbar_demux_001_src3_ready,         --            in.ready
			in_valid          => cmd_xbar_demux_001_src3_valid,         --              .valid
			in_startofpacket  => cmd_xbar_demux_001_src3_startofpacket, --              .startofpacket
			in_endofpacket    => cmd_xbar_demux_001_src3_endofpacket,   --              .endofpacket
			in_channel        => cmd_xbar_demux_001_src3_channel,       --              .channel
			in_data           => cmd_xbar_demux_001_src3_data,          --              .data
			out_ready         => crosser_out_ready,                     --           out.ready
			out_valid         => crosser_out_valid,                     --              .valid
			out_startofpacket => crosser_out_startofpacket,             --              .startofpacket
			out_endofpacket   => crosser_out_endofpacket,               --              .endofpacket
			out_channel       => crosser_out_channel,                   --              .channel
			out_data          => crosser_out_data,                      --              .data
			in_empty          => '0',                                   --   (terminated)
			in_error          => '0',                                   --   (terminated)
			out_empty         => open,                                  --   (terminated)
			out_error         => open                                   --   (terminated)
		);

	crosser_001 : component altera_avalon_st_handshake_clock_crosser
		generic map (
			DATA_WIDTH          => 104,
			BITS_PER_SYMBOL     => 104,
			USE_PACKETS         => 1,
			USE_CHANNEL         => 1,
			CHANNEL_WIDTH       => 33,
			USE_ERROR           => 0,
			ERROR_WIDTH         => 1,
			VALID_SYNC_DEPTH    => 2,
			READY_SYNC_DEPTH    => 2,
			USE_OUTPUT_PIPELINE => 0
		)
		port map (
			in_clk            => clk_50_clk,                            --        in_clk.clk
			in_reset          => rst_controller_001_reset_out_reset,    --  in_clk_reset.reset
			out_clk           => pll_c0_clk,                            --       out_clk.clk
			out_reset         => rst_controller_reset_out_reset,        -- out_clk_reset.reset
			in_ready          => rsp_xbar_demux_003_src0_ready,         --            in.ready
			in_valid          => rsp_xbar_demux_003_src0_valid,         --              .valid
			in_startofpacket  => rsp_xbar_demux_003_src0_startofpacket, --              .startofpacket
			in_endofpacket    => rsp_xbar_demux_003_src0_endofpacket,   --              .endofpacket
			in_channel        => rsp_xbar_demux_003_src0_channel,       --              .channel
			in_data           => rsp_xbar_demux_003_src0_data,          --              .data
			out_ready         => crosser_001_out_ready,                 --           out.ready
			out_valid         => crosser_001_out_valid,                 --              .valid
			out_startofpacket => crosser_001_out_startofpacket,         --              .startofpacket
			out_endofpacket   => crosser_001_out_endofpacket,           --              .endofpacket
			out_channel       => crosser_001_out_channel,               --              .channel
			out_data          => crosser_001_out_data,                  --              .data
			in_empty          => '0',                                   --   (terminated)
			in_error          => '0',                                   --   (terminated)
			out_empty         => open,                                  --   (terminated)
			out_error         => open                                   --   (terminated)
		);

	irq_mapper : component NIOSIImicro_irq_mapper
		port map (
			clk            => pll_c0_clk,                     --        clk.clk
			reset          => rst_controller_reset_out_reset, --  clk_reset.reset
			receiver0_irq  => irq_mapper_receiver0_irq,       --  receiver0.irq
			receiver1_irq  => irq_mapper_receiver1_irq,       --  receiver1.irq
			receiver2_irq  => irq_mapper_receiver2_irq,       --  receiver2.irq
			receiver3_irq  => irq_mapper_receiver3_irq,       --  receiver3.irq
			receiver4_irq  => irq_mapper_receiver4_irq,       --  receiver4.irq
			receiver5_irq  => irq_mapper_receiver5_irq,       --  receiver5.irq
			receiver6_irq  => irq_mapper_receiver6_irq,       --  receiver6.irq
			receiver7_irq  => irq_mapper_receiver7_irq,       --  receiver7.irq
			receiver8_irq  => irq_mapper_receiver8_irq,       --  receiver8.irq
			receiver9_irq  => irq_mapper_receiver9_irq,       --  receiver9.irq
			receiver10_irq => irq_mapper_receiver10_irq,      -- receiver10.irq
			receiver11_irq => irq_mapper_receiver11_irq,      -- receiver11.irq
			receiver12_irq => irq_mapper_receiver12_irq,      -- receiver12.irq
			receiver13_irq => irq_mapper_receiver13_irq,      -- receiver13.irq
			receiver14_irq => irq_mapper_receiver14_irq,      -- receiver14.irq
			receiver15_irq => irq_mapper_receiver15_irq,      -- receiver15.irq
			sender_irq     => cpu_d_irq_irq                   --     sender.irq
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	sdram_s1_translator_avalon_anti_slave_0_write_ports_inv <= not sdram_s1_translator_avalon_anti_slave_0_write;

	sdram_s1_translator_avalon_anti_slave_0_read_ports_inv <= not sdram_s1_translator_avalon_anti_slave_0_read;

	sdram_s1_translator_avalon_anti_slave_0_byteenable_ports_inv <= not sdram_s1_translator_avalon_anti_slave_0_byteenable;

	uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv <= not timer_0_s1_translator_avalon_anti_slave_0_write;

	timer_1_s1_translator_avalon_anti_slave_0_write_ports_inv <= not timer_1_s1_translator_avalon_anti_slave_0_write;

	pio_in_key_edge_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_in_key_edge_s1_translator_avalon_anti_slave_0_write;

	pio_in_ext_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_in_ext_s1_translator_avalon_anti_slave_0_write;

	pio_out_red_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_out_red_s1_translator_avalon_anti_slave_0_write;

	pio_out_green_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_out_green_s1_translator_avalon_anti_slave_0_write;

	pio_out_ext_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_out_ext_s1_translator_avalon_anti_slave_0_write;

	pio_async_reset_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_async_reset_s1_translator_avalon_anti_slave_0_write;

	pio_en_mux_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_en_mux_s1_translator_avalon_anti_slave_0_write;

	pio_direc_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_direc_s1_translator_avalon_anti_slave_0_write;

	pio_direc_ram_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_direc_ram_s1_translator_avalon_anti_slave_0_write;

	pio_wr_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_wr_s1_translator_avalon_anti_slave_0_write;

	pio_sel_salida_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_sel_salida_s1_translator_avalon_anti_slave_0_write;

	pio_datos_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_datos_s1_translator_avalon_anti_slave_0_write;

	pio_compara_int_0_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_compara_int_0_s1_translator_avalon_anti_slave_0_write;

	pio_compara_int_1_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_compara_int_1_s1_translator_avalon_anti_slave_0_write;

	pio_compara_int_2_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_compara_int_2_s1_translator_avalon_anti_slave_0_write;

	pio_compara_int_3_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_compara_int_3_s1_translator_avalon_anti_slave_0_write;

	pio_compara_int_4_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_compara_int_4_s1_translator_avalon_anti_slave_0_write;

	pio_captura_0_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_captura_0_s1_translator_avalon_anti_slave_0_write;

	pio_captura_1_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_captura_1_s1_translator_avalon_anti_slave_0_write;

	pio_captura_2_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_captura_2_s1_translator_avalon_anti_slave_0_write;

	pio_captura_3_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_captura_3_s1_translator_avalon_anti_slave_0_write;

	pio_captura_4_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_captura_4_s1_translator_avalon_anti_slave_0_write;

	pio_in_32_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_in_32_s1_translator_avalon_anti_slave_0_write;

	dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect_ports_inv <= not dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;

	dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write_ports_inv <= not dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write;

	dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read_ports_inv <= not dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of NIOSIImicro
